module registers(
  input        clk,
  input        rst,
  input        we,
  input  [7:0] dataw,
  input  [6:0] addr,
  output [7:0] datar,
  input  [3:0] regr_0,
  output [7:0] regwr_0,
  output [7:0] regwr_1,
  output [7:0] regwr_2,
  output [7:0] regwr_3,
  output [7:0] regwr_4,
  output [7:0] regwr_5,
  output [7:0] regwr_6,
  output [7:0] regwr_7,
  output [7:0] regwr_8,
  output [7:0] regwr_9,
  output [7:0] regwr_10,
  output [7:0] regwr_11,
  output [7:0] regwr_12,
  output [7:0] regwr_13,
  output [7:0] regwr_14,
  output [7:0] regwr_15,
  output [7:0] regwr_16,
  output [7:0] regwr_17,
  output [7:0] regwr_18,
  output [7:0] regwr_19,
  output [7:0] regwr_20,
  output [7:0] regwr_21,
  output [7:0] regwr_22,
  output [7:0] regwr_23,
  output [7:0] regwr_24,
  output [7:0] regwr_25,
  output [7:0] regwr_26,
  output [7:0] regwr_27,
  output [7:0] regwr_28,
  output [7:0] regwr_29,
  output [7:0] regwr_30,
  output [7:0] regwr_31,
  output [7:0] regwr_32,
  output [7:0] regwr_33,
  output [7:0] regwr_34,
  output [7:0] regwr_35,
  output [7:0] regwr_36,
  output [7:0] regwr_37,
  output [7:0] regwr_38,
  output [7:0] regwr_39,
  output [7:0] regwr_40,
  output [7:0] regwr_41,
  output [7:0] regwr_42,
  output [7:0] regwr_43,
  output [7:0] regwr_44,
  output [7:0] regwr_45,
  output [7:0] regwr_46,
  output [7:0] regwr_47,
  output [7:0] regwr_48,
  output [7:0] regwr_49,
  output [7:0] regwr_50,
  output [7:0] regwr_51,
  output [7:0] regwr_52,
  output [7:0] regwr_53,
  output [7:0] regwr_54,
  output [7:0] regwr_55,
  output [7:0] regwr_56,
  output [7:0] regwr_57,
  output [7:0] regwr_58,
  output [7:0] regwr_59,
  output [7:0] regwr_60,
  output [7:0] regwr_61,
  output [7:0] regwr_62,
  output [7:0] regwr_63,
  output [7:0] regwr_64,
  output [7:0] regwr_65,
  output [7:0] regwr_66,
  output [7:0] regwr_67,
  output [7:0] regwr_68,
  output [7:0] regwr_69,
  output [7:0] regwr_70,
  output [7:0] regwr_71,
  output [7:0] regwr_72,
  output [7:0] regwr_73,
  output [7:0] regwr_74,
  output [7:0] regwr_75,
  output [7:0] regwr_76,
  output [7:0] regwr_77,
  output [7:0] regwr_78,
  output [7:0] regwr_79,
  output [7:0] regwr_80,
  output [7:0] regwr_81,
  output [7:0] regwr_82,
  output [7:0] regwr_83,
  output [7:0] regwr_84,
  output [7:0] regwr_85,
  output [7:0] regwr_86,
  output [7:0] regwr_87,
  output [7:0] regwr_88,
  output [7:0] regwr_89,
  output [7:0] regwr_90,
  output [7:0] regwr_91,
  output [7:0] regwr_92,
  output [7:0] regwr_93,
  output [7:0] regwr_94,
  output [7:0] regwr_95,
  output [7:0] regwr_96,
  output [7:0] regwr_97,
  output [7:0] regwr_98,
  output [7:0] regwr_99,
  output [7:0] regwr_100,
  output [7:0] regwr_101,
  output [7:0] regwr_102,
  output [7:0] regwr_103,
  output [7:0] regwr_104,
  output [7:0] regwr_105,
  output [7:0] regwr_106,
  output [7:0] regwr_107,
  output [7:0] regwr_108,
  output [7:0] regwr_109,
  output [7:0] regwr_110,
  output [7:0] regwr_111,
  output [7:0] regwr_112,
  output [7:0] regwr_113,
  output [7:0] regwr_114,
  output [7:0] regwr_115,
  output [7:0] regwr_116,
  output [7:0] regwr_117,
  output [7:0] regwr_118,
  output [7:0] regwr_119,
  output [7:0] regwr_120
);
  reg [7:0] _T; // @[registers.scala 40:43]
  reg [31:0] _RAND_0;
  wire  _T_1 = addr == 7'h0; // @[registers.scala 41:39]
  wire  _T_2 = we & _T_1; // @[registers.scala 41:33]
  reg [7:0] _T_3; // @[registers.scala 40:43]
  reg [31:0] _RAND_1;
  wire  _T_4 = addr == 7'h1; // @[registers.scala 41:39]
  wire  _T_5 = we & _T_4; // @[registers.scala 41:33]
  reg [7:0] _T_6; // @[registers.scala 40:43]
  reg [31:0] _RAND_2;
  wire  _T_7 = addr == 7'h2; // @[registers.scala 41:39]
  wire  _T_8 = we & _T_7; // @[registers.scala 41:33]
  reg [7:0] _T_9; // @[registers.scala 40:43]
  reg [31:0] _RAND_3;
  wire  _T_10 = addr == 7'h3; // @[registers.scala 41:39]
  wire  _T_11 = we & _T_10; // @[registers.scala 41:33]
  reg [7:0] _T_12; // @[registers.scala 40:43]
  reg [31:0] _RAND_4;
  wire  _T_13 = addr == 7'h4; // @[registers.scala 41:39]
  wire  _T_14 = we & _T_13; // @[registers.scala 41:33]
  reg [7:0] _T_15; // @[registers.scala 40:43]
  reg [31:0] _RAND_5;
  wire  _T_16 = addr == 7'h5; // @[registers.scala 41:39]
  wire  _T_17 = we & _T_16; // @[registers.scala 41:33]
  reg [7:0] _T_18; // @[registers.scala 40:43]
  reg [31:0] _RAND_6;
  wire  _T_19 = addr == 7'h6; // @[registers.scala 41:39]
  wire  _T_20 = we & _T_19; // @[registers.scala 41:33]
  reg [7:0] _T_21; // @[registers.scala 40:43]
  reg [31:0] _RAND_7;
  wire  _T_22 = addr == 7'h7; // @[registers.scala 41:39]
  wire  _T_23 = we & _T_22; // @[registers.scala 41:33]
  reg [7:0] _T_24; // @[registers.scala 40:43]
  reg [31:0] _RAND_8;
  wire  _T_25 = addr == 7'h8; // @[registers.scala 41:39]
  wire  _T_26 = we & _T_25; // @[registers.scala 41:33]
  reg [7:0] _T_27; // @[registers.scala 40:43]
  reg [31:0] _RAND_9;
  wire  _T_28 = addr == 7'h9; // @[registers.scala 41:39]
  wire  _T_29 = we & _T_28; // @[registers.scala 41:33]
  reg [7:0] _T_30; // @[registers.scala 40:43]
  reg [31:0] _RAND_10;
  wire  _T_31 = addr == 7'ha; // @[registers.scala 41:39]
  wire  _T_32 = we & _T_31; // @[registers.scala 41:33]
  reg [7:0] _T_33; // @[registers.scala 40:43]
  reg [31:0] _RAND_11;
  wire  _T_34 = addr == 7'hb; // @[registers.scala 41:39]
  wire  _T_35 = we & _T_34; // @[registers.scala 41:33]
  reg [7:0] _T_36; // @[registers.scala 40:43]
  reg [31:0] _RAND_12;
  wire  _T_37 = addr == 7'hc; // @[registers.scala 41:39]
  wire  _T_38 = we & _T_37; // @[registers.scala 41:33]
  reg [7:0] _T_39; // @[registers.scala 40:43]
  reg [31:0] _RAND_13;
  wire  _T_40 = addr == 7'hd; // @[registers.scala 41:39]
  wire  _T_41 = we & _T_40; // @[registers.scala 41:33]
  reg [7:0] _T_42; // @[registers.scala 40:43]
  reg [31:0] _RAND_14;
  wire  _T_43 = addr == 7'he; // @[registers.scala 41:39]
  wire  _T_44 = we & _T_43; // @[registers.scala 41:33]
  reg [7:0] _T_45; // @[registers.scala 40:43]
  reg [31:0] _RAND_15;
  wire  _T_46 = addr == 7'hf; // @[registers.scala 41:39]
  wire  _T_47 = we & _T_46; // @[registers.scala 41:33]
  reg [7:0] _T_48; // @[registers.scala 40:43]
  reg [31:0] _RAND_16;
  wire  _T_49 = addr == 7'h10; // @[registers.scala 41:39]
  wire  _T_50 = we & _T_49; // @[registers.scala 41:33]
  reg [7:0] _T_51; // @[registers.scala 40:43]
  reg [31:0] _RAND_17;
  wire  _T_52 = addr == 7'h11; // @[registers.scala 41:39]
  wire  _T_53 = we & _T_52; // @[registers.scala 41:33]
  reg [7:0] _T_54; // @[registers.scala 40:43]
  reg [31:0] _RAND_18;
  wire  _T_55 = addr == 7'h12; // @[registers.scala 41:39]
  wire  _T_56 = we & _T_55; // @[registers.scala 41:33]
  reg [7:0] _T_57; // @[registers.scala 40:43]
  reg [31:0] _RAND_19;
  wire  _T_58 = addr == 7'h13; // @[registers.scala 41:39]
  wire  _T_59 = we & _T_58; // @[registers.scala 41:33]
  reg [7:0] _T_60; // @[registers.scala 40:43]
  reg [31:0] _RAND_20;
  wire  _T_61 = addr == 7'h14; // @[registers.scala 41:39]
  wire  _T_62 = we & _T_61; // @[registers.scala 41:33]
  reg [7:0] _T_63; // @[registers.scala 40:43]
  reg [31:0] _RAND_21;
  wire  _T_64 = addr == 7'h15; // @[registers.scala 41:39]
  wire  _T_65 = we & _T_64; // @[registers.scala 41:33]
  reg [7:0] _T_66; // @[registers.scala 40:43]
  reg [31:0] _RAND_22;
  wire  _T_67 = addr == 7'h16; // @[registers.scala 41:39]
  wire  _T_68 = we & _T_67; // @[registers.scala 41:33]
  reg [7:0] _T_69; // @[registers.scala 40:43]
  reg [31:0] _RAND_23;
  wire  _T_70 = addr == 7'h17; // @[registers.scala 41:39]
  wire  _T_71 = we & _T_70; // @[registers.scala 41:33]
  reg [7:0] _T_72; // @[registers.scala 40:43]
  reg [31:0] _RAND_24;
  wire  _T_73 = addr == 7'h18; // @[registers.scala 41:39]
  wire  _T_74 = we & _T_73; // @[registers.scala 41:33]
  reg [7:0] _T_75; // @[registers.scala 40:43]
  reg [31:0] _RAND_25;
  wire  _T_76 = addr == 7'h19; // @[registers.scala 41:39]
  wire  _T_77 = we & _T_76; // @[registers.scala 41:33]
  reg [7:0] _T_78; // @[registers.scala 40:43]
  reg [31:0] _RAND_26;
  wire  _T_79 = addr == 7'h1a; // @[registers.scala 41:39]
  wire  _T_80 = we & _T_79; // @[registers.scala 41:33]
  reg [7:0] _T_81; // @[registers.scala 40:43]
  reg [31:0] _RAND_27;
  wire  _T_82 = addr == 7'h1b; // @[registers.scala 41:39]
  wire  _T_83 = we & _T_82; // @[registers.scala 41:33]
  reg [7:0] _T_84; // @[registers.scala 40:43]
  reg [31:0] _RAND_28;
  wire  _T_85 = addr == 7'h1c; // @[registers.scala 41:39]
  wire  _T_86 = we & _T_85; // @[registers.scala 41:33]
  reg [7:0] _T_87; // @[registers.scala 40:43]
  reg [31:0] _RAND_29;
  wire  _T_88 = addr == 7'h1d; // @[registers.scala 41:39]
  wire  _T_89 = we & _T_88; // @[registers.scala 41:33]
  reg [7:0] _T_90; // @[registers.scala 40:43]
  reg [31:0] _RAND_30;
  wire  _T_91 = addr == 7'h1e; // @[registers.scala 41:39]
  wire  _T_92 = we & _T_91; // @[registers.scala 41:33]
  reg [7:0] _T_93; // @[registers.scala 40:43]
  reg [31:0] _RAND_31;
  wire  _T_94 = addr == 7'h1f; // @[registers.scala 41:39]
  wire  _T_95 = we & _T_94; // @[registers.scala 41:33]
  reg [7:0] _T_96; // @[registers.scala 40:43]
  reg [31:0] _RAND_32;
  wire  _T_97 = addr == 7'h20; // @[registers.scala 41:39]
  wire  _T_98 = we & _T_97; // @[registers.scala 41:33]
  reg [7:0] _T_99; // @[registers.scala 40:43]
  reg [31:0] _RAND_33;
  wire  _T_100 = addr == 7'h21; // @[registers.scala 41:39]
  wire  _T_101 = we & _T_100; // @[registers.scala 41:33]
  reg [7:0] _T_102; // @[registers.scala 40:43]
  reg [31:0] _RAND_34;
  wire  _T_103 = addr == 7'h22; // @[registers.scala 41:39]
  wire  _T_104 = we & _T_103; // @[registers.scala 41:33]
  reg [7:0] _T_105; // @[registers.scala 40:43]
  reg [31:0] _RAND_35;
  wire  _T_106 = addr == 7'h23; // @[registers.scala 41:39]
  wire  _T_107 = we & _T_106; // @[registers.scala 41:33]
  reg [7:0] _T_108; // @[registers.scala 40:43]
  reg [31:0] _RAND_36;
  wire  _T_109 = addr == 7'h24; // @[registers.scala 41:39]
  wire  _T_110 = we & _T_109; // @[registers.scala 41:33]
  reg [7:0] _T_111; // @[registers.scala 40:43]
  reg [31:0] _RAND_37;
  wire  _T_112 = addr == 7'h25; // @[registers.scala 41:39]
  wire  _T_113 = we & _T_112; // @[registers.scala 41:33]
  reg [7:0] _T_114; // @[registers.scala 40:43]
  reg [31:0] _RAND_38;
  wire  _T_115 = addr == 7'h26; // @[registers.scala 41:39]
  wire  _T_116 = we & _T_115; // @[registers.scala 41:33]
  reg [7:0] _T_117; // @[registers.scala 40:43]
  reg [31:0] _RAND_39;
  wire  _T_118 = addr == 7'h27; // @[registers.scala 41:39]
  wire  _T_119 = we & _T_118; // @[registers.scala 41:33]
  reg [7:0] _T_120; // @[registers.scala 40:43]
  reg [31:0] _RAND_40;
  wire  _T_121 = addr == 7'h28; // @[registers.scala 41:39]
  wire  _T_122 = we & _T_121; // @[registers.scala 41:33]
  reg [7:0] _T_123; // @[registers.scala 40:43]
  reg [31:0] _RAND_41;
  wire  _T_124 = addr == 7'h29; // @[registers.scala 41:39]
  wire  _T_125 = we & _T_124; // @[registers.scala 41:33]
  reg [7:0] _T_126; // @[registers.scala 40:43]
  reg [31:0] _RAND_42;
  wire  _T_127 = addr == 7'h2a; // @[registers.scala 41:39]
  wire  _T_128 = we & _T_127; // @[registers.scala 41:33]
  reg [7:0] _T_129; // @[registers.scala 40:43]
  reg [31:0] _RAND_43;
  wire  _T_130 = addr == 7'h2b; // @[registers.scala 41:39]
  wire  _T_131 = we & _T_130; // @[registers.scala 41:33]
  reg [7:0] _T_132; // @[registers.scala 40:43]
  reg [31:0] _RAND_44;
  wire  _T_133 = addr == 7'h2c; // @[registers.scala 41:39]
  wire  _T_134 = we & _T_133; // @[registers.scala 41:33]
  reg [7:0] _T_135; // @[registers.scala 40:43]
  reg [31:0] _RAND_45;
  wire  _T_136 = addr == 7'h2d; // @[registers.scala 41:39]
  wire  _T_137 = we & _T_136; // @[registers.scala 41:33]
  reg [7:0] _T_138; // @[registers.scala 40:43]
  reg [31:0] _RAND_46;
  wire  _T_139 = addr == 7'h2e; // @[registers.scala 41:39]
  wire  _T_140 = we & _T_139; // @[registers.scala 41:33]
  reg [7:0] _T_141; // @[registers.scala 40:43]
  reg [31:0] _RAND_47;
  wire  _T_142 = addr == 7'h2f; // @[registers.scala 41:39]
  wire  _T_143 = we & _T_142; // @[registers.scala 41:33]
  reg [7:0] _T_144; // @[registers.scala 40:43]
  reg [31:0] _RAND_48;
  wire  _T_145 = addr == 7'h30; // @[registers.scala 41:39]
  wire  _T_146 = we & _T_145; // @[registers.scala 41:33]
  reg [7:0] _T_147; // @[registers.scala 40:43]
  reg [31:0] _RAND_49;
  wire  _T_148 = addr == 7'h31; // @[registers.scala 41:39]
  wire  _T_149 = we & _T_148; // @[registers.scala 41:33]
  reg [7:0] _T_150; // @[registers.scala 40:43]
  reg [31:0] _RAND_50;
  wire  _T_151 = addr == 7'h32; // @[registers.scala 41:39]
  wire  _T_152 = we & _T_151; // @[registers.scala 41:33]
  reg [7:0] _T_153; // @[registers.scala 40:43]
  reg [31:0] _RAND_51;
  wire  _T_154 = addr == 7'h33; // @[registers.scala 41:39]
  wire  _T_155 = we & _T_154; // @[registers.scala 41:33]
  reg [7:0] _T_156; // @[registers.scala 40:43]
  reg [31:0] _RAND_52;
  wire  _T_157 = addr == 7'h34; // @[registers.scala 41:39]
  wire  _T_158 = we & _T_157; // @[registers.scala 41:33]
  reg [7:0] _T_159; // @[registers.scala 40:43]
  reg [31:0] _RAND_53;
  wire  _T_160 = addr == 7'h35; // @[registers.scala 41:39]
  wire  _T_161 = we & _T_160; // @[registers.scala 41:33]
  reg [7:0] _T_162; // @[registers.scala 40:43]
  reg [31:0] _RAND_54;
  wire  _T_163 = addr == 7'h36; // @[registers.scala 41:39]
  wire  _T_164 = we & _T_163; // @[registers.scala 41:33]
  reg [7:0] _T_165; // @[registers.scala 40:43]
  reg [31:0] _RAND_55;
  wire  _T_166 = addr == 7'h37; // @[registers.scala 41:39]
  wire  _T_167 = we & _T_166; // @[registers.scala 41:33]
  reg [7:0] _T_168; // @[registers.scala 40:43]
  reg [31:0] _RAND_56;
  wire  _T_169 = addr == 7'h38; // @[registers.scala 41:39]
  wire  _T_170 = we & _T_169; // @[registers.scala 41:33]
  reg [7:0] _T_171; // @[registers.scala 40:43]
  reg [31:0] _RAND_57;
  wire  _T_172 = addr == 7'h39; // @[registers.scala 41:39]
  wire  _T_173 = we & _T_172; // @[registers.scala 41:33]
  reg [7:0] _T_174; // @[registers.scala 40:43]
  reg [31:0] _RAND_58;
  wire  _T_175 = addr == 7'h3a; // @[registers.scala 41:39]
  wire  _T_176 = we & _T_175; // @[registers.scala 41:33]
  reg [7:0] _T_177; // @[registers.scala 40:43]
  reg [31:0] _RAND_59;
  wire  _T_178 = addr == 7'h3b; // @[registers.scala 41:39]
  wire  _T_179 = we & _T_178; // @[registers.scala 41:33]
  reg [7:0] _T_180; // @[registers.scala 40:43]
  reg [31:0] _RAND_60;
  wire  _T_181 = addr == 7'h3c; // @[registers.scala 41:39]
  wire  _T_182 = we & _T_181; // @[registers.scala 41:33]
  reg [7:0] _T_183; // @[registers.scala 40:43]
  reg [31:0] _RAND_61;
  wire  _T_184 = addr == 7'h3d; // @[registers.scala 41:39]
  wire  _T_185 = we & _T_184; // @[registers.scala 41:33]
  reg [7:0] _T_186; // @[registers.scala 40:43]
  reg [31:0] _RAND_62;
  wire  _T_187 = addr == 7'h3e; // @[registers.scala 41:39]
  wire  _T_188 = we & _T_187; // @[registers.scala 41:33]
  reg [7:0] _T_189; // @[registers.scala 40:43]
  reg [31:0] _RAND_63;
  wire  _T_190 = addr == 7'h3f; // @[registers.scala 41:39]
  wire  _T_191 = we & _T_190; // @[registers.scala 41:33]
  reg [7:0] _T_192; // @[registers.scala 40:43]
  reg [31:0] _RAND_64;
  wire  _T_193 = addr == 7'h40; // @[registers.scala 41:39]
  wire  _T_194 = we & _T_193; // @[registers.scala 41:33]
  reg [7:0] _T_195; // @[registers.scala 40:43]
  reg [31:0] _RAND_65;
  wire  _T_196 = addr == 7'h41; // @[registers.scala 41:39]
  wire  _T_197 = we & _T_196; // @[registers.scala 41:33]
  reg [7:0] _T_198; // @[registers.scala 40:43]
  reg [31:0] _RAND_66;
  wire  _T_199 = addr == 7'h42; // @[registers.scala 41:39]
  wire  _T_200 = we & _T_199; // @[registers.scala 41:33]
  reg [7:0] _T_201; // @[registers.scala 40:43]
  reg [31:0] _RAND_67;
  wire  _T_202 = addr == 7'h43; // @[registers.scala 41:39]
  wire  _T_203 = we & _T_202; // @[registers.scala 41:33]
  reg [7:0] _T_204; // @[registers.scala 40:43]
  reg [31:0] _RAND_68;
  wire  _T_205 = addr == 7'h44; // @[registers.scala 41:39]
  wire  _T_206 = we & _T_205; // @[registers.scala 41:33]
  reg [7:0] _T_207; // @[registers.scala 40:43]
  reg [31:0] _RAND_69;
  wire  _T_208 = addr == 7'h45; // @[registers.scala 41:39]
  wire  _T_209 = we & _T_208; // @[registers.scala 41:33]
  reg [7:0] _T_210; // @[registers.scala 40:43]
  reg [31:0] _RAND_70;
  wire  _T_211 = addr == 7'h46; // @[registers.scala 41:39]
  wire  _T_212 = we & _T_211; // @[registers.scala 41:33]
  reg [7:0] _T_213; // @[registers.scala 40:43]
  reg [31:0] _RAND_71;
  wire  _T_214 = addr == 7'h47; // @[registers.scala 41:39]
  wire  _T_215 = we & _T_214; // @[registers.scala 41:33]
  reg [7:0] _T_216; // @[registers.scala 40:43]
  reg [31:0] _RAND_72;
  wire  _T_217 = addr == 7'h48; // @[registers.scala 41:39]
  wire  _T_218 = we & _T_217; // @[registers.scala 41:33]
  reg [7:0] _T_219; // @[registers.scala 40:43]
  reg [31:0] _RAND_73;
  wire  _T_220 = addr == 7'h49; // @[registers.scala 41:39]
  wire  _T_221 = we & _T_220; // @[registers.scala 41:33]
  reg [7:0] _T_222; // @[registers.scala 40:43]
  reg [31:0] _RAND_74;
  wire  _T_223 = addr == 7'h4a; // @[registers.scala 41:39]
  wire  _T_224 = we & _T_223; // @[registers.scala 41:33]
  reg [7:0] _T_225; // @[registers.scala 40:43]
  reg [31:0] _RAND_75;
  wire  _T_226 = addr == 7'h4b; // @[registers.scala 41:39]
  wire  _T_227 = we & _T_226; // @[registers.scala 41:33]
  reg [7:0] _T_228; // @[registers.scala 40:43]
  reg [31:0] _RAND_76;
  wire  _T_229 = addr == 7'h4c; // @[registers.scala 41:39]
  wire  _T_230 = we & _T_229; // @[registers.scala 41:33]
  reg [7:0] _T_231; // @[registers.scala 40:43]
  reg [31:0] _RAND_77;
  wire  _T_232 = addr == 7'h4d; // @[registers.scala 41:39]
  wire  _T_233 = we & _T_232; // @[registers.scala 41:33]
  reg [7:0] _T_234; // @[registers.scala 40:43]
  reg [31:0] _RAND_78;
  wire  _T_235 = addr == 7'h4e; // @[registers.scala 41:39]
  wire  _T_236 = we & _T_235; // @[registers.scala 41:33]
  reg [7:0] _T_237; // @[registers.scala 40:43]
  reg [31:0] _RAND_79;
  wire  _T_238 = addr == 7'h4f; // @[registers.scala 41:39]
  wire  _T_239 = we & _T_238; // @[registers.scala 41:33]
  reg [7:0] _T_240; // @[registers.scala 40:43]
  reg [31:0] _RAND_80;
  wire  _T_241 = addr == 7'h50; // @[registers.scala 41:39]
  wire  _T_242 = we & _T_241; // @[registers.scala 41:33]
  reg [7:0] _T_243; // @[registers.scala 40:43]
  reg [31:0] _RAND_81;
  wire  _T_244 = addr == 7'h51; // @[registers.scala 41:39]
  wire  _T_245 = we & _T_244; // @[registers.scala 41:33]
  reg [7:0] _T_246; // @[registers.scala 40:43]
  reg [31:0] _RAND_82;
  wire  _T_247 = addr == 7'h52; // @[registers.scala 41:39]
  wire  _T_248 = we & _T_247; // @[registers.scala 41:33]
  reg [7:0] _T_249; // @[registers.scala 40:43]
  reg [31:0] _RAND_83;
  wire  _T_250 = addr == 7'h53; // @[registers.scala 41:39]
  wire  _T_251 = we & _T_250; // @[registers.scala 41:33]
  reg [7:0] _T_252; // @[registers.scala 40:43]
  reg [31:0] _RAND_84;
  wire  _T_253 = addr == 7'h54; // @[registers.scala 41:39]
  wire  _T_254 = we & _T_253; // @[registers.scala 41:33]
  reg [7:0] _T_255; // @[registers.scala 40:43]
  reg [31:0] _RAND_85;
  wire  _T_256 = addr == 7'h55; // @[registers.scala 41:39]
  wire  _T_257 = we & _T_256; // @[registers.scala 41:33]
  reg [7:0] _T_258; // @[registers.scala 40:43]
  reg [31:0] _RAND_86;
  wire  _T_259 = addr == 7'h56; // @[registers.scala 41:39]
  wire  _T_260 = we & _T_259; // @[registers.scala 41:33]
  reg [7:0] _T_261; // @[registers.scala 40:43]
  reg [31:0] _RAND_87;
  wire  _T_262 = addr == 7'h57; // @[registers.scala 41:39]
  wire  _T_263 = we & _T_262; // @[registers.scala 41:33]
  reg [7:0] _T_264; // @[registers.scala 40:43]
  reg [31:0] _RAND_88;
  wire  _T_265 = addr == 7'h58; // @[registers.scala 41:39]
  wire  _T_266 = we & _T_265; // @[registers.scala 41:33]
  reg [7:0] _T_267; // @[registers.scala 40:43]
  reg [31:0] _RAND_89;
  wire  _T_268 = addr == 7'h59; // @[registers.scala 41:39]
  wire  _T_269 = we & _T_268; // @[registers.scala 41:33]
  reg [7:0] _T_270; // @[registers.scala 40:43]
  reg [31:0] _RAND_90;
  wire  _T_271 = addr == 7'h5a; // @[registers.scala 41:39]
  wire  _T_272 = we & _T_271; // @[registers.scala 41:33]
  reg [7:0] _T_273; // @[registers.scala 40:43]
  reg [31:0] _RAND_91;
  wire  _T_274 = addr == 7'h5b; // @[registers.scala 41:39]
  wire  _T_275 = we & _T_274; // @[registers.scala 41:33]
  reg [7:0] _T_276; // @[registers.scala 40:43]
  reg [31:0] _RAND_92;
  wire  _T_277 = addr == 7'h5c; // @[registers.scala 41:39]
  wire  _T_278 = we & _T_277; // @[registers.scala 41:33]
  reg [7:0] _T_279; // @[registers.scala 40:43]
  reg [31:0] _RAND_93;
  wire  _T_280 = addr == 7'h5d; // @[registers.scala 41:39]
  wire  _T_281 = we & _T_280; // @[registers.scala 41:33]
  reg [7:0] _T_282; // @[registers.scala 40:43]
  reg [31:0] _RAND_94;
  wire  _T_283 = addr == 7'h5e; // @[registers.scala 41:39]
  wire  _T_284 = we & _T_283; // @[registers.scala 41:33]
  reg [7:0] _T_285; // @[registers.scala 40:43]
  reg [31:0] _RAND_95;
  wire  _T_286 = addr == 7'h5f; // @[registers.scala 41:39]
  wire  _T_287 = we & _T_286; // @[registers.scala 41:33]
  reg [7:0] _T_288; // @[registers.scala 40:43]
  reg [31:0] _RAND_96;
  wire  _T_289 = addr == 7'h60; // @[registers.scala 41:39]
  wire  _T_290 = we & _T_289; // @[registers.scala 41:33]
  reg [7:0] _T_291; // @[registers.scala 40:43]
  reg [31:0] _RAND_97;
  wire  _T_292 = addr == 7'h61; // @[registers.scala 41:39]
  wire  _T_293 = we & _T_292; // @[registers.scala 41:33]
  reg [7:0] _T_294; // @[registers.scala 40:43]
  reg [31:0] _RAND_98;
  wire  _T_295 = addr == 7'h62; // @[registers.scala 41:39]
  wire  _T_296 = we & _T_295; // @[registers.scala 41:33]
  reg [7:0] _T_297; // @[registers.scala 40:43]
  reg [31:0] _RAND_99;
  wire  _T_298 = addr == 7'h63; // @[registers.scala 41:39]
  wire  _T_299 = we & _T_298; // @[registers.scala 41:33]
  reg [7:0] _T_300; // @[registers.scala 40:43]
  reg [31:0] _RAND_100;
  wire  _T_301 = addr == 7'h64; // @[registers.scala 41:39]
  wire  _T_302 = we & _T_301; // @[registers.scala 41:33]
  reg [7:0] _T_303; // @[registers.scala 40:43]
  reg [31:0] _RAND_101;
  wire  _T_304 = addr == 7'h65; // @[registers.scala 41:39]
  wire  _T_305 = we & _T_304; // @[registers.scala 41:33]
  reg [7:0] _T_306; // @[registers.scala 40:43]
  reg [31:0] _RAND_102;
  wire  _T_307 = addr == 7'h66; // @[registers.scala 41:39]
  wire  _T_308 = we & _T_307; // @[registers.scala 41:33]
  reg [7:0] _T_309; // @[registers.scala 40:43]
  reg [31:0] _RAND_103;
  wire  _T_310 = addr == 7'h67; // @[registers.scala 41:39]
  wire  _T_311 = we & _T_310; // @[registers.scala 41:33]
  reg [7:0] _T_312; // @[registers.scala 40:43]
  reg [31:0] _RAND_104;
  wire  _T_313 = addr == 7'h68; // @[registers.scala 41:39]
  wire  _T_314 = we & _T_313; // @[registers.scala 41:33]
  reg [7:0] _T_315; // @[registers.scala 40:43]
  reg [31:0] _RAND_105;
  wire  _T_316 = addr == 7'h69; // @[registers.scala 41:39]
  wire  _T_317 = we & _T_316; // @[registers.scala 41:33]
  reg [7:0] _T_318; // @[registers.scala 40:43]
  reg [31:0] _RAND_106;
  wire  _T_319 = addr == 7'h6a; // @[registers.scala 41:39]
  wire  _T_320 = we & _T_319; // @[registers.scala 41:33]
  reg [7:0] _T_321; // @[registers.scala 40:43]
  reg [31:0] _RAND_107;
  wire  _T_322 = addr == 7'h6b; // @[registers.scala 41:39]
  wire  _T_323 = we & _T_322; // @[registers.scala 41:33]
  reg [7:0] _T_324; // @[registers.scala 40:43]
  reg [31:0] _RAND_108;
  wire  _T_325 = addr == 7'h6c; // @[registers.scala 41:39]
  wire  _T_326 = we & _T_325; // @[registers.scala 41:33]
  reg [7:0] _T_327; // @[registers.scala 40:43]
  reg [31:0] _RAND_109;
  wire  _T_328 = addr == 7'h6d; // @[registers.scala 41:39]
  wire  _T_329 = we & _T_328; // @[registers.scala 41:33]
  reg [7:0] _T_330; // @[registers.scala 40:43]
  reg [31:0] _RAND_110;
  wire  _T_331 = addr == 7'h6e; // @[registers.scala 41:39]
  wire  _T_332 = we & _T_331; // @[registers.scala 41:33]
  reg [7:0] _T_333; // @[registers.scala 40:43]
  reg [31:0] _RAND_111;
  wire  _T_334 = addr == 7'h6f; // @[registers.scala 41:39]
  wire  _T_335 = we & _T_334; // @[registers.scala 41:33]
  reg [7:0] _T_336; // @[registers.scala 40:43]
  reg [31:0] _RAND_112;
  wire  _T_337 = addr == 7'h70; // @[registers.scala 41:39]
  wire  _T_338 = we & _T_337; // @[registers.scala 41:33]
  reg [7:0] _T_339; // @[registers.scala 40:43]
  reg [31:0] _RAND_113;
  wire  _T_340 = addr == 7'h71; // @[registers.scala 41:39]
  wire  _T_341 = we & _T_340; // @[registers.scala 41:33]
  reg [7:0] _T_342; // @[registers.scala 40:43]
  reg [31:0] _RAND_114;
  wire  _T_343 = addr == 7'h72; // @[registers.scala 41:39]
  wire  _T_344 = we & _T_343; // @[registers.scala 41:33]
  reg [7:0] _T_345; // @[registers.scala 40:43]
  reg [31:0] _RAND_115;
  wire  _T_346 = addr == 7'h73; // @[registers.scala 41:39]
  wire  _T_347 = we & _T_346; // @[registers.scala 41:33]
  reg [7:0] _T_348; // @[registers.scala 40:43]
  reg [31:0] _RAND_116;
  wire  _T_349 = addr == 7'h74; // @[registers.scala 41:39]
  wire  _T_350 = we & _T_349; // @[registers.scala 41:33]
  reg [7:0] _T_351; // @[registers.scala 40:43]
  reg [31:0] _RAND_117;
  wire  _T_352 = addr == 7'h75; // @[registers.scala 41:39]
  wire  _T_353 = we & _T_352; // @[registers.scala 41:33]
  reg [7:0] _T_354; // @[registers.scala 40:43]
  reg [31:0] _RAND_118;
  wire  _T_355 = addr == 7'h76; // @[registers.scala 41:39]
  wire  _T_356 = we & _T_355; // @[registers.scala 41:33]
  reg [7:0] _T_357; // @[registers.scala 40:43]
  reg [31:0] _RAND_119;
  wire  _T_358 = addr == 7'h77; // @[registers.scala 41:39]
  wire  _T_359 = we & _T_358; // @[registers.scala 41:33]
  reg [7:0] _T_360; // @[registers.scala 40:43]
  reg [31:0] _RAND_120;
  wire  _T_361 = addr == 7'h78; // @[registers.scala 41:39]
  wire  _T_362 = we & _T_361; // @[registers.scala 41:33]
  reg [7:0] _T_365_0; // @[registers.scala 51:39]
  reg [31:0] _RAND_121;
  wire [55:0] _T_372 = {_T_18,_T_15,_T_12,_T_9,_T_6,_T_3,_T}; // @[registers.scala 61:68]
  wire [119:0] _T_380 = {_T_42,_T_39,_T_36,_T_33,_T_30,_T_27,_T_24,_T_21,_T_372}; // @[registers.scala 61:68]
  wire [55:0] _T_386 = {_T_63,_T_60,_T_57,_T_54,_T_51,_T_48,_T_45}; // @[registers.scala 61:68]
  wire [239:0] _T_395 = {_T_87,_T_84,_T_81,_T_78,_T_75,_T_72,_T_69,_T_66,_T_386,_T_380}; // @[registers.scala 61:68]
  wire [55:0] _T_401 = {_T_108,_T_105,_T_102,_T_99,_T_96,_T_93,_T_90}; // @[registers.scala 61:68]
  wire [119:0] _T_409 = {_T_132,_T_129,_T_126,_T_123,_T_120,_T_117,_T_114,_T_111,_T_401}; // @[registers.scala 61:68]
  wire [55:0] _T_415 = {_T_153,_T_150,_T_147,_T_144,_T_141,_T_138,_T_135}; // @[registers.scala 61:68]
  wire [239:0] _T_424 = {_T_177,_T_174,_T_171,_T_168,_T_165,_T_162,_T_159,_T_156,_T_415,_T_409}; // @[registers.scala 61:68]
  wire [55:0] _T_431 = {_T_198,_T_195,_T_192,_T_189,_T_186,_T_183,_T_180}; // @[registers.scala 61:68]
  wire [119:0] _T_439 = {_T_222,_T_219,_T_216,_T_213,_T_210,_T_207,_T_204,_T_201,_T_431}; // @[registers.scala 61:68]
  wire [55:0] _T_445 = {_T_243,_T_240,_T_237,_T_234,_T_231,_T_228,_T_225}; // @[registers.scala 61:68]
  wire [239:0] _T_454 = {_T_267,_T_264,_T_261,_T_258,_T_255,_T_252,_T_249,_T_246,_T_445,_T_439}; // @[registers.scala 61:68]
  wire [55:0] _T_460 = {_T_288,_T_285,_T_282,_T_279,_T_276,_T_273,_T_270}; // @[registers.scala 61:68]
  wire [119:0] _T_468 = {_T_312,_T_309,_T_306,_T_303,_T_300,_T_297,_T_294,_T_291,_T_460}; // @[registers.scala 61:68]
  wire [63:0] _T_475 = {_T_336,_T_333,_T_330,_T_327,_T_324,_T_321,_T_318,_T_315}; // @[registers.scala 61:68]
  wire [247:0] _T_484 = {_T_360,_T_357,_T_354,_T_351,_T_348,_T_345,_T_342,_T_339,_T_475,_T_468}; // @[registers.scala 61:68]
  wire [975:0] _T_487 = {_T_365_0,_T_484,_T_454,_T_424,_T_395}; // @[Cat.scala 30:58]
  reg [7:0] _T_612; // @[registers.scala 63:37]
  reg [31:0] _RAND_122;
  assign datar = _T_612; // @[registers.scala 64:22]
  assign regwr_0 = _T; // @[registers.scala 46:33]
  assign regwr_1 = _T_3; // @[registers.scala 46:33]
  assign regwr_2 = _T_6; // @[registers.scala 46:33]
  assign regwr_3 = _T_9; // @[registers.scala 46:33]
  assign regwr_4 = _T_12; // @[registers.scala 46:33]
  assign regwr_5 = _T_15; // @[registers.scala 46:33]
  assign regwr_6 = _T_18; // @[registers.scala 46:33]
  assign regwr_7 = _T_21; // @[registers.scala 46:33]
  assign regwr_8 = _T_24; // @[registers.scala 46:33]
  assign regwr_9 = _T_27; // @[registers.scala 46:33]
  assign regwr_10 = _T_30; // @[registers.scala 46:33]
  assign regwr_11 = _T_33; // @[registers.scala 46:33]
  assign regwr_12 = _T_36; // @[registers.scala 46:33]
  assign regwr_13 = _T_39; // @[registers.scala 46:33]
  assign regwr_14 = _T_42; // @[registers.scala 46:33]
  assign regwr_15 = _T_45; // @[registers.scala 46:33]
  assign regwr_16 = _T_48; // @[registers.scala 46:33]
  assign regwr_17 = _T_51; // @[registers.scala 46:33]
  assign regwr_18 = _T_54; // @[registers.scala 46:33]
  assign regwr_19 = _T_57; // @[registers.scala 46:33]
  assign regwr_20 = _T_60; // @[registers.scala 46:33]
  assign regwr_21 = _T_63; // @[registers.scala 46:33]
  assign regwr_22 = _T_66; // @[registers.scala 46:33]
  assign regwr_23 = _T_69; // @[registers.scala 46:33]
  assign regwr_24 = _T_72; // @[registers.scala 46:33]
  assign regwr_25 = _T_75; // @[registers.scala 46:33]
  assign regwr_26 = _T_78; // @[registers.scala 46:33]
  assign regwr_27 = _T_81; // @[registers.scala 46:33]
  assign regwr_28 = _T_84; // @[registers.scala 46:33]
  assign regwr_29 = _T_87; // @[registers.scala 46:33]
  assign regwr_30 = _T_90; // @[registers.scala 46:33]
  assign regwr_31 = _T_93; // @[registers.scala 46:33]
  assign regwr_32 = _T_96; // @[registers.scala 46:33]
  assign regwr_33 = _T_99; // @[registers.scala 46:33]
  assign regwr_34 = _T_102; // @[registers.scala 46:33]
  assign regwr_35 = _T_105; // @[registers.scala 46:33]
  assign regwr_36 = _T_108; // @[registers.scala 46:33]
  assign regwr_37 = _T_111; // @[registers.scala 46:33]
  assign regwr_38 = _T_114; // @[registers.scala 46:33]
  assign regwr_39 = _T_117; // @[registers.scala 46:33]
  assign regwr_40 = _T_120; // @[registers.scala 46:33]
  assign regwr_41 = _T_123; // @[registers.scala 46:33]
  assign regwr_42 = _T_126; // @[registers.scala 46:33]
  assign regwr_43 = _T_129; // @[registers.scala 46:33]
  assign regwr_44 = _T_132; // @[registers.scala 46:33]
  assign regwr_45 = _T_135; // @[registers.scala 46:33]
  assign regwr_46 = _T_138; // @[registers.scala 46:33]
  assign regwr_47 = _T_141; // @[registers.scala 46:33]
  assign regwr_48 = _T_144; // @[registers.scala 46:33]
  assign regwr_49 = _T_147; // @[registers.scala 46:33]
  assign regwr_50 = _T_150; // @[registers.scala 46:33]
  assign regwr_51 = _T_153; // @[registers.scala 46:33]
  assign regwr_52 = _T_156; // @[registers.scala 46:33]
  assign regwr_53 = _T_159; // @[registers.scala 46:33]
  assign regwr_54 = _T_162; // @[registers.scala 46:33]
  assign regwr_55 = _T_165; // @[registers.scala 46:33]
  assign regwr_56 = _T_168; // @[registers.scala 46:33]
  assign regwr_57 = _T_171; // @[registers.scala 46:33]
  assign regwr_58 = _T_174; // @[registers.scala 46:33]
  assign regwr_59 = _T_177; // @[registers.scala 46:33]
  assign regwr_60 = _T_180; // @[registers.scala 46:33]
  assign regwr_61 = _T_183; // @[registers.scala 46:33]
  assign regwr_62 = _T_186; // @[registers.scala 46:33]
  assign regwr_63 = _T_189; // @[registers.scala 46:33]
  assign regwr_64 = _T_192; // @[registers.scala 46:33]
  assign regwr_65 = _T_195; // @[registers.scala 46:33]
  assign regwr_66 = _T_198; // @[registers.scala 46:33]
  assign regwr_67 = _T_201; // @[registers.scala 46:33]
  assign regwr_68 = _T_204; // @[registers.scala 46:33]
  assign regwr_69 = _T_207; // @[registers.scala 46:33]
  assign regwr_70 = _T_210; // @[registers.scala 46:33]
  assign regwr_71 = _T_213; // @[registers.scala 46:33]
  assign regwr_72 = _T_216; // @[registers.scala 46:33]
  assign regwr_73 = _T_219; // @[registers.scala 46:33]
  assign regwr_74 = _T_222; // @[registers.scala 46:33]
  assign regwr_75 = _T_225; // @[registers.scala 46:33]
  assign regwr_76 = _T_228; // @[registers.scala 46:33]
  assign regwr_77 = _T_231; // @[registers.scala 46:33]
  assign regwr_78 = _T_234; // @[registers.scala 46:33]
  assign regwr_79 = _T_237; // @[registers.scala 46:33]
  assign regwr_80 = _T_240; // @[registers.scala 46:33]
  assign regwr_81 = _T_243; // @[registers.scala 46:33]
  assign regwr_82 = _T_246; // @[registers.scala 46:33]
  assign regwr_83 = _T_249; // @[registers.scala 46:33]
  assign regwr_84 = _T_252; // @[registers.scala 46:33]
  assign regwr_85 = _T_255; // @[registers.scala 46:33]
  assign regwr_86 = _T_258; // @[registers.scala 46:33]
  assign regwr_87 = _T_261; // @[registers.scala 46:33]
  assign regwr_88 = _T_264; // @[registers.scala 46:33]
  assign regwr_89 = _T_267; // @[registers.scala 46:33]
  assign regwr_90 = _T_270; // @[registers.scala 46:33]
  assign regwr_91 = _T_273; // @[registers.scala 46:33]
  assign regwr_92 = _T_276; // @[registers.scala 46:33]
  assign regwr_93 = _T_279; // @[registers.scala 46:33]
  assign regwr_94 = _T_282; // @[registers.scala 46:33]
  assign regwr_95 = _T_285; // @[registers.scala 46:33]
  assign regwr_96 = _T_288; // @[registers.scala 46:33]
  assign regwr_97 = _T_291; // @[registers.scala 46:33]
  assign regwr_98 = _T_294; // @[registers.scala 46:33]
  assign regwr_99 = _T_297; // @[registers.scala 46:33]
  assign regwr_100 = _T_300; // @[registers.scala 46:33]
  assign regwr_101 = _T_303; // @[registers.scala 46:33]
  assign regwr_102 = _T_306; // @[registers.scala 46:33]
  assign regwr_103 = _T_309; // @[registers.scala 46:33]
  assign regwr_104 = _T_312; // @[registers.scala 46:33]
  assign regwr_105 = _T_315; // @[registers.scala 46:33]
  assign regwr_106 = _T_318; // @[registers.scala 46:33]
  assign regwr_107 = _T_321; // @[registers.scala 46:33]
  assign regwr_108 = _T_324; // @[registers.scala 46:33]
  assign regwr_109 = _T_327; // @[registers.scala 46:33]
  assign regwr_110 = _T_330; // @[registers.scala 46:33]
  assign regwr_111 = _T_333; // @[registers.scala 46:33]
  assign regwr_112 = _T_336; // @[registers.scala 46:33]
  assign regwr_113 = _T_339; // @[registers.scala 46:33]
  assign regwr_114 = _T_342; // @[registers.scala 46:33]
  assign regwr_115 = _T_345; // @[registers.scala 46:33]
  assign regwr_116 = _T_348; // @[registers.scala 46:33]
  assign regwr_117 = _T_351; // @[registers.scala 46:33]
  assign regwr_118 = _T_354; // @[registers.scala 46:33]
  assign regwr_119 = _T_357; // @[registers.scala 46:33]
  assign regwr_120 = _T_360; // @[registers.scala 46:33]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_3 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_6 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_9 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_12 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_15 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_18 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_21 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_24 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_27 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_30 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_33 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_36 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_39 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_42 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_45 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_48 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_51 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_54 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_57 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_60 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_63 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_66 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_69 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_72 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_75 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_78 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_81 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_84 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_87 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_90 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_93 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_96 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_99 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_102 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_105 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_108 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_111 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_114 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_117 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_120 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_123 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_126 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_129 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_132 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_135 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_138 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_141 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_144 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_147 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_150 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_153 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_156 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_159 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_162 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_165 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_168 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_171 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_174 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_177 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_180 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_183 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_186 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_189 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_192 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_195 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_198 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_201 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_204 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_207 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_210 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_213 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_216 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_219 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_222 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_225 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_228 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_231 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_234 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_237 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_240 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_243 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_246 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_249 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_252 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_255 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_258 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_261 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_264 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_267 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_270 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_273 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_276 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_279 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_282 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_285 = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_288 = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_291 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_294 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_297 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_300 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_303 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_306 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_309 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_312 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_315 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_318 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_321 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_324 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_327 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_330 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_333 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_336 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_339 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_342 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_345 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_348 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_351 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_354 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_357 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_360 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_365_0 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_612 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  if (rst) begin
    _T = 8'h0;
  end
  if (rst) begin
    _T_3 = 8'h0;
  end
  if (rst) begin
    _T_6 = 8'h0;
  end
  if (rst) begin
    _T_9 = 8'h0;
  end
  if (rst) begin
    _T_12 = 8'h0;
  end
  if (rst) begin
    _T_15 = 8'h0;
  end
  if (rst) begin
    _T_18 = 8'h0;
  end
  if (rst) begin
    _T_21 = 8'h0;
  end
  if (rst) begin
    _T_24 = 8'h0;
  end
  if (rst) begin
    _T_27 = 8'h0;
  end
  if (rst) begin
    _T_30 = 8'h0;
  end
  if (rst) begin
    _T_33 = 8'h0;
  end
  if (rst) begin
    _T_36 = 8'h0;
  end
  if (rst) begin
    _T_39 = 8'h0;
  end
  if (rst) begin
    _T_42 = 8'h0;
  end
  if (rst) begin
    _T_45 = 8'h0;
  end
  if (rst) begin
    _T_48 = 8'h0;
  end
  if (rst) begin
    _T_51 = 8'h0;
  end
  if (rst) begin
    _T_54 = 8'h0;
  end
  if (rst) begin
    _T_57 = 8'h0;
  end
  if (rst) begin
    _T_60 = 8'h0;
  end
  if (rst) begin
    _T_63 = 8'h0;
  end
  if (rst) begin
    _T_66 = 8'h0;
  end
  if (rst) begin
    _T_69 = 8'h0;
  end
  if (rst) begin
    _T_72 = 8'h0;
  end
  if (rst) begin
    _T_75 = 8'h0;
  end
  if (rst) begin
    _T_78 = 8'h0;
  end
  if (rst) begin
    _T_81 = 8'h0;
  end
  if (rst) begin
    _T_84 = 8'h0;
  end
  if (rst) begin
    _T_87 = 8'h0;
  end
  if (rst) begin
    _T_90 = 8'h0;
  end
  if (rst) begin
    _T_93 = 8'h0;
  end
  if (rst) begin
    _T_96 = 8'h0;
  end
  if (rst) begin
    _T_99 = 8'h0;
  end
  if (rst) begin
    _T_102 = 8'h0;
  end
  if (rst) begin
    _T_105 = 8'h0;
  end
  if (rst) begin
    _T_108 = 8'h0;
  end
  if (rst) begin
    _T_111 = 8'h0;
  end
  if (rst) begin
    _T_114 = 8'h0;
  end
  if (rst) begin
    _T_117 = 8'h0;
  end
  if (rst) begin
    _T_120 = 8'h0;
  end
  if (rst) begin
    _T_123 = 8'h0;
  end
  if (rst) begin
    _T_126 = 8'h0;
  end
  if (rst) begin
    _T_129 = 8'h0;
  end
  if (rst) begin
    _T_132 = 8'h0;
  end
  if (rst) begin
    _T_135 = 8'h0;
  end
  if (rst) begin
    _T_138 = 8'h0;
  end
  if (rst) begin
    _T_141 = 8'h0;
  end
  if (rst) begin
    _T_144 = 8'h0;
  end
  if (rst) begin
    _T_147 = 8'h0;
  end
  if (rst) begin
    _T_150 = 8'h0;
  end
  if (rst) begin
    _T_153 = 8'h0;
  end
  if (rst) begin
    _T_156 = 8'h0;
  end
  if (rst) begin
    _T_159 = 8'h0;
  end
  if (rst) begin
    _T_162 = 8'h0;
  end
  if (rst) begin
    _T_165 = 8'h0;
  end
  if (rst) begin
    _T_168 = 8'h0;
  end
  if (rst) begin
    _T_171 = 8'h0;
  end
  if (rst) begin
    _T_174 = 8'h0;
  end
  if (rst) begin
    _T_177 = 8'h0;
  end
  if (rst) begin
    _T_180 = 8'h0;
  end
  if (rst) begin
    _T_183 = 8'h0;
  end
  if (rst) begin
    _T_186 = 8'h0;
  end
  if (rst) begin
    _T_189 = 8'h0;
  end
  if (rst) begin
    _T_192 = 8'h0;
  end
  if (rst) begin
    _T_195 = 8'h0;
  end
  if (rst) begin
    _T_198 = 8'h0;
  end
  if (rst) begin
    _T_201 = 8'h0;
  end
  if (rst) begin
    _T_204 = 8'h0;
  end
  if (rst) begin
    _T_207 = 8'h0;
  end
  if (rst) begin
    _T_210 = 8'h0;
  end
  if (rst) begin
    _T_213 = 8'h0;
  end
  if (rst) begin
    _T_216 = 8'h0;
  end
  if (rst) begin
    _T_219 = 8'h0;
  end
  if (rst) begin
    _T_222 = 8'h0;
  end
  if (rst) begin
    _T_225 = 8'h0;
  end
  if (rst) begin
    _T_228 = 8'h0;
  end
  if (rst) begin
    _T_231 = 8'h0;
  end
  if (rst) begin
    _T_234 = 8'h0;
  end
  if (rst) begin
    _T_237 = 8'h0;
  end
  if (rst) begin
    _T_240 = 8'h0;
  end
  if (rst) begin
    _T_243 = 8'h0;
  end
  if (rst) begin
    _T_246 = 8'h0;
  end
  if (rst) begin
    _T_249 = 8'h0;
  end
  if (rst) begin
    _T_252 = 8'h0;
  end
  if (rst) begin
    _T_255 = 8'h0;
  end
  if (rst) begin
    _T_258 = 8'h0;
  end
  if (rst) begin
    _T_261 = 8'h0;
  end
  if (rst) begin
    _T_264 = 8'h0;
  end
  if (rst) begin
    _T_267 = 8'h0;
  end
  if (rst) begin
    _T_270 = 8'h0;
  end
  if (rst) begin
    _T_273 = 8'h0;
  end
  if (rst) begin
    _T_276 = 8'h0;
  end
  if (rst) begin
    _T_279 = 8'h0;
  end
  if (rst) begin
    _T_282 = 8'h0;
  end
  if (rst) begin
    _T_285 = 8'h0;
  end
  if (rst) begin
    _T_288 = 8'h0;
  end
  if (rst) begin
    _T_291 = 8'h0;
  end
  if (rst) begin
    _T_294 = 8'h0;
  end
  if (rst) begin
    _T_297 = 8'h0;
  end
  if (rst) begin
    _T_300 = 8'h0;
  end
  if (rst) begin
    _T_303 = 8'h0;
  end
  if (rst) begin
    _T_306 = 8'h0;
  end
  if (rst) begin
    _T_309 = 8'h0;
  end
  if (rst) begin
    _T_312 = 8'h0;
  end
  if (rst) begin
    _T_315 = 8'h0;
  end
  if (rst) begin
    _T_318 = 8'h0;
  end
  if (rst) begin
    _T_321 = 8'h0;
  end
  if (rst) begin
    _T_324 = 8'h0;
  end
  if (rst) begin
    _T_327 = 8'h0;
  end
  if (rst) begin
    _T_330 = 8'h0;
  end
  if (rst) begin
    _T_333 = 8'h0;
  end
  if (rst) begin
    _T_336 = 8'h0;
  end
  if (rst) begin
    _T_339 = 8'h0;
  end
  if (rst) begin
    _T_342 = 8'h0;
  end
  if (rst) begin
    _T_345 = 8'h0;
  end
  if (rst) begin
    _T_348 = 8'h0;
  end
  if (rst) begin
    _T_351 = 8'h0;
  end
  if (rst) begin
    _T_354 = 8'h0;
  end
  if (rst) begin
    _T_357 = 8'h0;
  end
  if (rst) begin
    _T_360 = 8'h0;
  end
  if (rst) begin
    _T_365_0 = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clk) begin
    if (7'h79 == addr) begin
      _T_612 <= _T_487[975:968];
    end else if (7'h78 == addr) begin
      _T_612 <= _T_487[967:960];
    end else if (7'h77 == addr) begin
      _T_612 <= _T_487[959:952];
    end else if (7'h76 == addr) begin
      _T_612 <= _T_487[951:944];
    end else if (7'h75 == addr) begin
      _T_612 <= _T_487[943:936];
    end else if (7'h74 == addr) begin
      _T_612 <= _T_487[935:928];
    end else if (7'h73 == addr) begin
      _T_612 <= _T_487[927:920];
    end else if (7'h72 == addr) begin
      _T_612 <= _T_487[919:912];
    end else if (7'h71 == addr) begin
      _T_612 <= _T_487[911:904];
    end else if (7'h70 == addr) begin
      _T_612 <= _T_487[903:896];
    end else if (7'h6f == addr) begin
      _T_612 <= _T_487[895:888];
    end else if (7'h6e == addr) begin
      _T_612 <= _T_487[887:880];
    end else if (7'h6d == addr) begin
      _T_612 <= _T_487[879:872];
    end else if (7'h6c == addr) begin
      _T_612 <= _T_487[871:864];
    end else if (7'h6b == addr) begin
      _T_612 <= _T_487[863:856];
    end else if (7'h6a == addr) begin
      _T_612 <= _T_487[855:848];
    end else if (7'h69 == addr) begin
      _T_612 <= _T_487[847:840];
    end else if (7'h68 == addr) begin
      _T_612 <= _T_487[839:832];
    end else if (7'h67 == addr) begin
      _T_612 <= _T_487[831:824];
    end else if (7'h66 == addr) begin
      _T_612 <= _T_487[823:816];
    end else if (7'h65 == addr) begin
      _T_612 <= _T_487[815:808];
    end else if (7'h64 == addr) begin
      _T_612 <= _T_487[807:800];
    end else if (7'h63 == addr) begin
      _T_612 <= _T_487[799:792];
    end else if (7'h62 == addr) begin
      _T_612 <= _T_487[791:784];
    end else if (7'h61 == addr) begin
      _T_612 <= _T_487[783:776];
    end else if (7'h60 == addr) begin
      _T_612 <= _T_487[775:768];
    end else if (7'h5f == addr) begin
      _T_612 <= _T_487[767:760];
    end else if (7'h5e == addr) begin
      _T_612 <= _T_487[759:752];
    end else if (7'h5d == addr) begin
      _T_612 <= _T_487[751:744];
    end else if (7'h5c == addr) begin
      _T_612 <= _T_487[743:736];
    end else if (7'h5b == addr) begin
      _T_612 <= _T_487[735:728];
    end else if (7'h5a == addr) begin
      _T_612 <= _T_487[727:720];
    end else if (7'h59 == addr) begin
      _T_612 <= _T_487[719:712];
    end else if (7'h58 == addr) begin
      _T_612 <= _T_487[711:704];
    end else if (7'h57 == addr) begin
      _T_612 <= _T_487[703:696];
    end else if (7'h56 == addr) begin
      _T_612 <= _T_487[695:688];
    end else if (7'h55 == addr) begin
      _T_612 <= _T_487[687:680];
    end else if (7'h54 == addr) begin
      _T_612 <= _T_487[679:672];
    end else if (7'h53 == addr) begin
      _T_612 <= _T_487[671:664];
    end else if (7'h52 == addr) begin
      _T_612 <= _T_487[663:656];
    end else if (7'h51 == addr) begin
      _T_612 <= _T_487[655:648];
    end else if (7'h50 == addr) begin
      _T_612 <= _T_487[647:640];
    end else if (7'h4f == addr) begin
      _T_612 <= _T_487[639:632];
    end else if (7'h4e == addr) begin
      _T_612 <= _T_487[631:624];
    end else if (7'h4d == addr) begin
      _T_612 <= _T_487[623:616];
    end else if (7'h4c == addr) begin
      _T_612 <= _T_487[615:608];
    end else if (7'h4b == addr) begin
      _T_612 <= _T_487[607:600];
    end else if (7'h4a == addr) begin
      _T_612 <= _T_487[599:592];
    end else if (7'h49 == addr) begin
      _T_612 <= _T_487[591:584];
    end else if (7'h48 == addr) begin
      _T_612 <= _T_487[583:576];
    end else if (7'h47 == addr) begin
      _T_612 <= _T_487[575:568];
    end else if (7'h46 == addr) begin
      _T_612 <= _T_487[567:560];
    end else if (7'h45 == addr) begin
      _T_612 <= _T_487[559:552];
    end else if (7'h44 == addr) begin
      _T_612 <= _T_487[551:544];
    end else if (7'h43 == addr) begin
      _T_612 <= _T_487[543:536];
    end else if (7'h42 == addr) begin
      _T_612 <= _T_487[535:528];
    end else if (7'h41 == addr) begin
      _T_612 <= _T_487[527:520];
    end else if (7'h40 == addr) begin
      _T_612 <= _T_487[519:512];
    end else if (7'h3f == addr) begin
      _T_612 <= _T_487[511:504];
    end else if (7'h3e == addr) begin
      _T_612 <= _T_487[503:496];
    end else if (7'h3d == addr) begin
      _T_612 <= _T_487[495:488];
    end else if (7'h3c == addr) begin
      _T_612 <= _T_487[487:480];
    end else if (7'h3b == addr) begin
      _T_612 <= _T_487[479:472];
    end else if (7'h3a == addr) begin
      _T_612 <= _T_487[471:464];
    end else if (7'h39 == addr) begin
      _T_612 <= _T_487[463:456];
    end else if (7'h38 == addr) begin
      _T_612 <= _T_487[455:448];
    end else if (7'h37 == addr) begin
      _T_612 <= _T_487[447:440];
    end else if (7'h36 == addr) begin
      _T_612 <= _T_487[439:432];
    end else if (7'h35 == addr) begin
      _T_612 <= _T_487[431:424];
    end else if (7'h34 == addr) begin
      _T_612 <= _T_487[423:416];
    end else if (7'h33 == addr) begin
      _T_612 <= _T_487[415:408];
    end else if (7'h32 == addr) begin
      _T_612 <= _T_487[407:400];
    end else if (7'h31 == addr) begin
      _T_612 <= _T_487[399:392];
    end else if (7'h30 == addr) begin
      _T_612 <= _T_487[391:384];
    end else if (7'h2f == addr) begin
      _T_612 <= _T_487[383:376];
    end else if (7'h2e == addr) begin
      _T_612 <= _T_487[375:368];
    end else if (7'h2d == addr) begin
      _T_612 <= _T_487[367:360];
    end else if (7'h2c == addr) begin
      _T_612 <= _T_487[359:352];
    end else if (7'h2b == addr) begin
      _T_612 <= _T_487[351:344];
    end else if (7'h2a == addr) begin
      _T_612 <= _T_487[343:336];
    end else if (7'h29 == addr) begin
      _T_612 <= _T_487[335:328];
    end else if (7'h28 == addr) begin
      _T_612 <= _T_487[327:320];
    end else if (7'h27 == addr) begin
      _T_612 <= _T_487[319:312];
    end else if (7'h26 == addr) begin
      _T_612 <= _T_487[311:304];
    end else if (7'h25 == addr) begin
      _T_612 <= _T_487[303:296];
    end else if (7'h24 == addr) begin
      _T_612 <= _T_487[295:288];
    end else if (7'h23 == addr) begin
      _T_612 <= _T_487[287:280];
    end else if (7'h22 == addr) begin
      _T_612 <= _T_487[279:272];
    end else if (7'h21 == addr) begin
      _T_612 <= _T_487[271:264];
    end else if (7'h20 == addr) begin
      _T_612 <= _T_487[263:256];
    end else if (7'h1f == addr) begin
      _T_612 <= _T_487[255:248];
    end else if (7'h1e == addr) begin
      _T_612 <= _T_487[247:240];
    end else if (7'h1d == addr) begin
      _T_612 <= _T_487[239:232];
    end else if (7'h1c == addr) begin
      _T_612 <= _T_487[231:224];
    end else if (7'h1b == addr) begin
      _T_612 <= _T_487[223:216];
    end else if (7'h1a == addr) begin
      _T_612 <= _T_487[215:208];
    end else if (7'h19 == addr) begin
      _T_612 <= _T_487[207:200];
    end else if (7'h18 == addr) begin
      _T_612 <= _T_487[199:192];
    end else if (7'h17 == addr) begin
      _T_612 <= _T_487[191:184];
    end else if (7'h16 == addr) begin
      _T_612 <= _T_487[183:176];
    end else if (7'h15 == addr) begin
      _T_612 <= _T_487[175:168];
    end else if (7'h14 == addr) begin
      _T_612 <= _T_487[167:160];
    end else if (7'h13 == addr) begin
      _T_612 <= _T_487[159:152];
    end else if (7'h12 == addr) begin
      _T_612 <= _T_487[151:144];
    end else if (7'h11 == addr) begin
      _T_612 <= _T_487[143:136];
    end else if (7'h10 == addr) begin
      _T_612 <= _T_487[135:128];
    end else if (7'hf == addr) begin
      _T_612 <= _T_487[127:120];
    end else if (7'he == addr) begin
      _T_612 <= _T_487[119:112];
    end else if (7'hd == addr) begin
      _T_612 <= _T_487[111:104];
    end else if (7'hc == addr) begin
      _T_612 <= _T_487[103:96];
    end else if (7'hb == addr) begin
      _T_612 <= _T_487[95:88];
    end else if (7'ha == addr) begin
      _T_612 <= _T_487[87:80];
    end else if (7'h9 == addr) begin
      _T_612 <= _T_487[79:72];
    end else if (7'h8 == addr) begin
      _T_612 <= _T_487[71:64];
    end else if (7'h7 == addr) begin
      _T_612 <= _T_487[63:56];
    end else if (7'h6 == addr) begin
      _T_612 <= _T_487[55:48];
    end else if (7'h5 == addr) begin
      _T_612 <= _T_487[47:40];
    end else if (7'h4 == addr) begin
      _T_612 <= _T_487[39:32];
    end else if (7'h3 == addr) begin
      _T_612 <= _T_487[31:24];
    end else if (7'h2 == addr) begin
      _T_612 <= _T_487[23:16];
    end else if (7'h1 == addr) begin
      _T_612 <= _T_487[15:8];
    end else begin
      _T_612 <= _T_487[7:0];
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T <= 8'h0;
    end else if (_T_2) begin
      _T <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_3 <= 8'h0;
    end else if (_T_5) begin
      _T_3 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_6 <= 8'h0;
    end else if (_T_8) begin
      _T_6 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_9 <= 8'h0;
    end else if (_T_11) begin
      _T_9 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_12 <= 8'h0;
    end else if (_T_14) begin
      _T_12 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_15 <= 8'h0;
    end else if (_T_17) begin
      _T_15 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_18 <= 8'h0;
    end else if (_T_20) begin
      _T_18 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_21 <= 8'h0;
    end else if (_T_23) begin
      _T_21 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_24 <= 8'h0;
    end else if (_T_26) begin
      _T_24 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_27 <= 8'h0;
    end else if (_T_29) begin
      _T_27 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_30 <= 8'h0;
    end else if (_T_32) begin
      _T_30 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_33 <= 8'h0;
    end else if (_T_35) begin
      _T_33 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_36 <= 8'h0;
    end else if (_T_38) begin
      _T_36 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_39 <= 8'h0;
    end else if (_T_41) begin
      _T_39 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_42 <= 8'h0;
    end else if (_T_44) begin
      _T_42 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_45 <= 8'h0;
    end else if (_T_47) begin
      _T_45 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_48 <= 8'h0;
    end else if (_T_50) begin
      _T_48 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_51 <= 8'h0;
    end else if (_T_53) begin
      _T_51 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_54 <= 8'h0;
    end else if (_T_56) begin
      _T_54 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_57 <= 8'h0;
    end else if (_T_59) begin
      _T_57 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_60 <= 8'h0;
    end else if (_T_62) begin
      _T_60 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_63 <= 8'h0;
    end else if (_T_65) begin
      _T_63 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_66 <= 8'h0;
    end else if (_T_68) begin
      _T_66 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_69 <= 8'h0;
    end else if (_T_71) begin
      _T_69 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_72 <= 8'h0;
    end else if (_T_74) begin
      _T_72 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_75 <= 8'h0;
    end else if (_T_77) begin
      _T_75 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_78 <= 8'h0;
    end else if (_T_80) begin
      _T_78 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_81 <= 8'h0;
    end else if (_T_83) begin
      _T_81 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_84 <= 8'h0;
    end else if (_T_86) begin
      _T_84 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_87 <= 8'h0;
    end else if (_T_89) begin
      _T_87 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_90 <= 8'h0;
    end else if (_T_92) begin
      _T_90 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_93 <= 8'h0;
    end else if (_T_95) begin
      _T_93 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_96 <= 8'h0;
    end else if (_T_98) begin
      _T_96 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_99 <= 8'h0;
    end else if (_T_101) begin
      _T_99 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_102 <= 8'h0;
    end else if (_T_104) begin
      _T_102 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_105 <= 8'h0;
    end else if (_T_107) begin
      _T_105 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_108 <= 8'h0;
    end else if (_T_110) begin
      _T_108 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_111 <= 8'h0;
    end else if (_T_113) begin
      _T_111 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_114 <= 8'h0;
    end else if (_T_116) begin
      _T_114 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_117 <= 8'h0;
    end else if (_T_119) begin
      _T_117 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_120 <= 8'h0;
    end else if (_T_122) begin
      _T_120 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_123 <= 8'h0;
    end else if (_T_125) begin
      _T_123 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_126 <= 8'h0;
    end else if (_T_128) begin
      _T_126 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_129 <= 8'h0;
    end else if (_T_131) begin
      _T_129 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_132 <= 8'h0;
    end else if (_T_134) begin
      _T_132 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_135 <= 8'h0;
    end else if (_T_137) begin
      _T_135 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_138 <= 8'h0;
    end else if (_T_140) begin
      _T_138 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_141 <= 8'h0;
    end else if (_T_143) begin
      _T_141 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_144 <= 8'h0;
    end else if (_T_146) begin
      _T_144 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_147 <= 8'h0;
    end else if (_T_149) begin
      _T_147 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_150 <= 8'h0;
    end else if (_T_152) begin
      _T_150 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_153 <= 8'h0;
    end else if (_T_155) begin
      _T_153 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_156 <= 8'h0;
    end else if (_T_158) begin
      _T_156 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_159 <= 8'h0;
    end else if (_T_161) begin
      _T_159 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_162 <= 8'h0;
    end else if (_T_164) begin
      _T_162 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_165 <= 8'h0;
    end else if (_T_167) begin
      _T_165 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_168 <= 8'h0;
    end else if (_T_170) begin
      _T_168 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_171 <= 8'h0;
    end else if (_T_173) begin
      _T_171 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_174 <= 8'h0;
    end else if (_T_176) begin
      _T_174 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_177 <= 8'h0;
    end else if (_T_179) begin
      _T_177 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_180 <= 8'h0;
    end else if (_T_182) begin
      _T_180 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_183 <= 8'h0;
    end else if (_T_185) begin
      _T_183 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_186 <= 8'h0;
    end else if (_T_188) begin
      _T_186 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_189 <= 8'h0;
    end else if (_T_191) begin
      _T_189 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_192 <= 8'h0;
    end else if (_T_194) begin
      _T_192 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_195 <= 8'h0;
    end else if (_T_197) begin
      _T_195 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_198 <= 8'h0;
    end else if (_T_200) begin
      _T_198 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_201 <= 8'h0;
    end else if (_T_203) begin
      _T_201 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_204 <= 8'h0;
    end else if (_T_206) begin
      _T_204 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_207 <= 8'h0;
    end else if (_T_209) begin
      _T_207 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_210 <= 8'h0;
    end else if (_T_212) begin
      _T_210 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_213 <= 8'h0;
    end else if (_T_215) begin
      _T_213 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_216 <= 8'h0;
    end else if (_T_218) begin
      _T_216 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_219 <= 8'h0;
    end else if (_T_221) begin
      _T_219 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_222 <= 8'h0;
    end else if (_T_224) begin
      _T_222 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_225 <= 8'h0;
    end else if (_T_227) begin
      _T_225 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_228 <= 8'h0;
    end else if (_T_230) begin
      _T_228 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_231 <= 8'h0;
    end else if (_T_233) begin
      _T_231 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_234 <= 8'h0;
    end else if (_T_236) begin
      _T_234 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_237 <= 8'h0;
    end else if (_T_239) begin
      _T_237 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_240 <= 8'h0;
    end else if (_T_242) begin
      _T_240 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_243 <= 8'h0;
    end else if (_T_245) begin
      _T_243 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_246 <= 8'h0;
    end else if (_T_248) begin
      _T_246 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_249 <= 8'h0;
    end else if (_T_251) begin
      _T_249 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_252 <= 8'h0;
    end else if (_T_254) begin
      _T_252 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_255 <= 8'h0;
    end else if (_T_257) begin
      _T_255 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_258 <= 8'h0;
    end else if (_T_260) begin
      _T_258 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_261 <= 8'h0;
    end else if (_T_263) begin
      _T_261 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_264 <= 8'h0;
    end else if (_T_266) begin
      _T_264 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_267 <= 8'h0;
    end else if (_T_269) begin
      _T_267 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_270 <= 8'h0;
    end else if (_T_272) begin
      _T_270 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_273 <= 8'h0;
    end else if (_T_275) begin
      _T_273 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_276 <= 8'h0;
    end else if (_T_278) begin
      _T_276 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_279 <= 8'h0;
    end else if (_T_281) begin
      _T_279 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_282 <= 8'h0;
    end else if (_T_284) begin
      _T_282 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_285 <= 8'h0;
    end else if (_T_287) begin
      _T_285 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_288 <= 8'h0;
    end else if (_T_290) begin
      _T_288 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_291 <= 8'h0;
    end else if (_T_293) begin
      _T_291 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_294 <= 8'h0;
    end else if (_T_296) begin
      _T_294 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_297 <= 8'h0;
    end else if (_T_299) begin
      _T_297 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_300 <= 8'h0;
    end else if (_T_302) begin
      _T_300 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_303 <= 8'h0;
    end else if (_T_305) begin
      _T_303 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_306 <= 8'h0;
    end else if (_T_308) begin
      _T_306 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_309 <= 8'h0;
    end else if (_T_311) begin
      _T_309 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_312 <= 8'h0;
    end else if (_T_314) begin
      _T_312 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_315 <= 8'h0;
    end else if (_T_317) begin
      _T_315 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_318 <= 8'h0;
    end else if (_T_320) begin
      _T_318 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_321 <= 8'h0;
    end else if (_T_323) begin
      _T_321 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_324 <= 8'h0;
    end else if (_T_326) begin
      _T_324 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_327 <= 8'h0;
    end else if (_T_329) begin
      _T_327 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_330 <= 8'h0;
    end else if (_T_332) begin
      _T_330 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_333 <= 8'h0;
    end else if (_T_335) begin
      _T_333 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_336 <= 8'h0;
    end else if (_T_338) begin
      _T_336 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_339 <= 8'h0;
    end else if (_T_341) begin
      _T_339 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_342 <= 8'h0;
    end else if (_T_344) begin
      _T_342 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_345 <= 8'h0;
    end else if (_T_347) begin
      _T_345 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_348 <= 8'h0;
    end else if (_T_350) begin
      _T_348 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_351 <= 8'h0;
    end else if (_T_353) begin
      _T_351 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_354 <= 8'h0;
    end else if (_T_356) begin
      _T_354 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_357 <= 8'h0;
    end else if (_T_359) begin
      _T_357 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_360 <= 8'h0;
    end else if (_T_362) begin
      _T_360 <= dataw;
    end
  end
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      _T_365_0 <= 8'h0;
    end else begin
      _T_365_0 <= {{4'd0}, regr_0};
    end
  end
endmodule