`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Universidad Industrial de Santander
// Engineer: Edward Silva
// 
// Create Date: 07/07/2021 
// Design Name: Network
// Module Name: Top
// Project Name: Library development for A-Connect
// Target Devices: Implementation on FPGA 
// 
//////////////////////////////////////////////////////////////////////////////////


module Top#( parameter number_image = 121, parameter size_word = 8)(
  input [7:0] regwr_0,
  input [7:0] regwr_1,
  input [7:0] regwr_2,
  input [7:0] regwr_3,
  input [7:0] regwr_4,
  input [7:0] regwr_5,
  input [7:0] regwr_6,
  input [7:0] regwr_7,
  input [7:0] regwr_8,
  input [7:0] regwr_9,
  input [7:0] regwr_10,
  input [7:0] regwr_11,
  input [7:0] regwr_12,
  input [7:0] regwr_13,
  input [7:0] regwr_14,
  input [7:0] regwr_15,
  input [7:0] regwr_16,
  input [7:0] regwr_17,
  input [7:0] regwr_18,
  input [7:0] regwr_19,
  input [7:0] regwr_20,
  input [7:0] regwr_21,
  input [7:0] regwr_22,
  input [7:0] regwr_23,
  input [7:0] regwr_24,
  input [7:0] regwr_25,
  input [7:0] regwr_26,
  input [7:0] regwr_27,
  input [7:0] regwr_28,
  input [7:0] regwr_29,
  input [7:0] regwr_30,
  input [7:0] regwr_31,
  input [7:0] regwr_32,
  input [7:0] regwr_33,
  input [7:0] regwr_34,
  input [7:0] regwr_35,
  input [7:0] regwr_36,
  input [7:0] regwr_37,
  input [7:0] regwr_38,
  input [7:0] regwr_39,
  input [7:0] regwr_40,
  input [7:0] regwr_41,
  input [7:0] regwr_42,
  input [7:0] regwr_43,
  input [7:0] regwr_44,
  input [7:0] regwr_45,
  input [7:0] regwr_46,
  input [7:0] regwr_47,
  input [7:0] regwr_48,
  input [7:0] regwr_49,
  input [7:0] regwr_50,
  input [7:0] regwr_51,
  input [7:0] regwr_52,
  input [7:0] regwr_53,
  input [7:0] regwr_54,
  input [7:0] regwr_55,
  input [7:0] regwr_56,
  input [7:0] regwr_57,
  input [7:0] regwr_58,
  input [7:0] regwr_59,
  input [7:0] regwr_60,
  input [7:0] regwr_61,
  input [7:0] regwr_62,
  input [7:0] regwr_63,
  input [7:0] regwr_64,
  input [7:0] regwr_65,
  input [7:0] regwr_66,
  input [7:0] regwr_67,
  input [7:0] regwr_68,
  input [7:0] regwr_69,
  input [7:0] regwr_70,
  input [7:0] regwr_71,
  input [7:0] regwr_72,
  input [7:0] regwr_73,
  input [7:0] regwr_74,
  input [7:0] regwr_75,
  input [7:0] regwr_76,
  input [7:0] regwr_77,
  input [7:0] regwr_78,
  input [7:0] regwr_79,
  input [7:0] regwr_80,
  input [7:0] regwr_81,
  input [7:0] regwr_82,
  input [7:0] regwr_83,
  input [7:0] regwr_84,
  input [7:0] regwr_85,
  input [7:0] regwr_86,
  input [7:0] regwr_87,
  input [7:0] regwr_88,
  input [7:0] regwr_89,
  input [7:0] regwr_90,
  input [7:0] regwr_91,
  input [7:0] regwr_92,
  input [7:0] regwr_93,
  input [7:0] regwr_94,
  input [7:0] regwr_95,
  input [7:0] regwr_96,
  input [7:0] regwr_97,
  input [7:0] regwr_98,
  input [7:0] regwr_99,
  input [7:0] regwr_100,
  input [7:0] regwr_101,
  input [7:0] regwr_102,
  input [7:0] regwr_103,
  input [7:0] regwr_104,
  input [7:0] regwr_105,
  input [7:0] regwr_106,
  input [7:0] regwr_107,
  input [7:0] regwr_108,
  input [7:0] regwr_109,
  input [7:0] regwr_110,
  input [7:0] regwr_111,
  input [7:0] regwr_112,
  input [7:0] regwr_113,
  input [7:0] regwr_114,
  input [7:0] regwr_115,
  input [7:0] regwr_116,
  input [7:0] regwr_117,
  input [7:0] regwr_118,
  input [7:0] regwr_119,
  input [7:0] regwr_120,
  
  output [3:0] regr_0
  
  );
  
  
  //******* Prueba con red del paper *******
  localparam number_output1 = 60; 
  localparam number_out = 10;
  
    //******* Acomodando las imagenes de entrada *******
  reg [size_word*number_image-1:0] Image; //Requerida como entrada de modulo neuron.v
  reg [number_image-1:0] Weight [0:number_output1-1];
  reg [number_output1-1:0] Weight_out [0:number_out-1];
  
  wire [2*size_word*number_output1-1:0]out_aux;
  wire [4*size_word*number_out-1:0]out_aux_out;
  
  //wire [18*number_output1-1:0]out_aux;
  //wire [2*18*number_out-1:0]out_aux_out;
  
  //******************************************
  //reg [3:0] scaling [0:47];
  //reg signed [3:0] offset [0:47];
  
  
  always@(*) 
  begin
	//Acomodando en un vector los pixeles de la imagen
	Image[7:0] = regwr_0; 
	Image[15:8] = regwr_1; 
	Image[23:16] = regwr_2; 
	Image[31:24] = regwr_3; 
	Image[39:32] = regwr_4; 
	Image[47:40] = regwr_5; 
	Image[55:48] = regwr_6; 
	Image[63:56] = regwr_7; 
	Image[71:64] = regwr_8; 
	Image[79:72] = regwr_9; 
	Image[87:80] = regwr_10; 
	Image[95:88] = regwr_11; 
	Image[103:96] = regwr_12; 
	Image[111:104] = regwr_13; 
	Image[119:112] = regwr_14; 
	Image[127:120] = regwr_15; 
	Image[135:128] = regwr_16; 
	Image[143:136] = regwr_17; 
	Image[151:144] = regwr_18; 
	Image[159:152] = regwr_19; 
	Image[167:160] = regwr_20; 
	Image[175:168] = regwr_21; 
	Image[183:176] = regwr_22; 
	Image[191:184] = regwr_23; 
	Image[199:192] = regwr_24; 
	Image[207:200] = regwr_25; 
	Image[215:208] = regwr_26; 
	Image[223:216] = regwr_27; 
	Image[231:224] = regwr_28; 
	Image[239:232] = regwr_29; 
	Image[247:240] = regwr_30; 
	Image[255:248] = regwr_31; 
	Image[263:256] = regwr_32; 
	Image[271:264] = regwr_33; 
	Image[279:272] = regwr_34; 
	Image[287:280] = regwr_35; 
	Image[295:288] = regwr_36; 
	Image[303:296] = regwr_37; 
	Image[311:304] = regwr_38; 
	Image[319:312] = regwr_39; 
	Image[327:320] = regwr_40; 
	Image[335:328] = regwr_41; 
	Image[343:336] = regwr_42; 
	Image[351:344] = regwr_43; 
	Image[359:352] = regwr_44; 
	Image[367:360] = regwr_45; 
	Image[375:368] = regwr_46; 
	Image[383:376] = regwr_47; 
	Image[391:384] = regwr_48; 
	Image[399:392] = regwr_49; 
	Image[407:400] = regwr_50; 
	Image[415:408] = regwr_51; 
	Image[423:416] = regwr_52; 
	Image[431:424] = regwr_53; 
	Image[439:432] = regwr_54; 
	Image[447:440] = regwr_55; 
	Image[455:448] = regwr_56; 
	Image[463:456] = regwr_57; 
	Image[471:464] = regwr_58; 
	Image[479:472] = regwr_59; 
	Image[487:480] = regwr_60; 
	Image[495:488] = regwr_61; 
	Image[503:496] = regwr_62; 
	Image[511:504] = regwr_63; 
	Image[519:512] = regwr_64; 
	Image[527:520] = regwr_65; 
	Image[535:528] = regwr_66; 
	Image[543:536] = regwr_67; 
	Image[551:544] = regwr_68; 
	Image[559:552] = regwr_69; 
	Image[567:560] = regwr_70; 
	Image[575:568] = regwr_71; 
	Image[583:576] = regwr_72; 
	Image[591:584] = regwr_73; 
	Image[599:592] = regwr_74; 
	Image[607:600] = regwr_75; 
	Image[615:608] = regwr_76; 
	Image[623:616] = regwr_77; 
	Image[631:624] = regwr_78; 
	Image[639:632] = regwr_79; 
	Image[647:640] = regwr_80; 
	Image[655:648] = regwr_81; 
	Image[663:656] = regwr_82; 
	Image[671:664] = regwr_83; 
	Image[679:672] = regwr_84; 
	Image[687:680] = regwr_85; 
	Image[695:688] = regwr_86; 
	Image[703:696] = regwr_87; 
	Image[711:704] = regwr_88; 
	Image[719:712] = regwr_89; 
	Image[727:720] = regwr_90; 
	Image[735:728] = regwr_91; 
	Image[743:736] = regwr_92; 
	Image[751:744] = regwr_93; 
	Image[759:752] = regwr_94; 
	Image[767:760] = regwr_95; 
	Image[775:768] = regwr_96; 
	Image[783:776] = regwr_97; 
	Image[791:784] = regwr_98; 
	Image[799:792] = regwr_99; 
	Image[807:800] = regwr_100; 
	Image[815:808] = regwr_101; 
	Image[823:816] = regwr_102; 
	Image[831:824] = regwr_103; 
	Image[839:832] = regwr_104; 
	Image[847:840] = regwr_105; 
	Image[855:848] = regwr_106; 
	Image[863:856] = regwr_107; 
	Image[871:864] = regwr_108; 
	Image[879:872] = regwr_109; 
	Image[887:880] = regwr_110; 
	Image[895:888] = regwr_111; 
	Image[903:896] = regwr_112; 
	Image[911:904] = regwr_113; 
	Image[919:912] = regwr_114; 
	Image[927:920] = regwr_115; 
	Image[935:928] = regwr_116; 
	Image[943:936] = regwr_117; 
	Image[951:944] = regwr_118; 
	Image[959:952] = regwr_119; 
	Image[967:960] = regwr_120; 
 
	
	//****** Net for Implementation ****** New function reshape Image
	 //Loading weight [60,121] : [output,input] with BatchNormalization
	 //****** Prueba con red del paper ******
	//Loading weight [60,121] : [output,input]
	Weight[0] = 121'b1010101010111001000100110110110110000010111010011001010000011111111100011000000010000011100110000000001110001101111110101;
	Weight[1] = 121'b1100001000111101111000101111111000000101100010000011110000010111011011101000101011000111111110010111011110000100001101010;
	Weight[2] = 121'b0001101010110001100001001011100000101011100101110001001100100110001000000001010011110000100011010101000111101110000111100;
	Weight[3] = 121'b1110000110001111111110100000000010010100011000000111111110011101101010000100001111111000000111000011001000001011100001010;
	Weight[4] = 121'b0100000000111100001101101011001100111110111111000101000100010000100111011111011000010100100000011000011100000001111010101;
	Weight[5] = 121'b1000110111010010110011010111110100001001111000111101111001100001101011100001100001000011110111110001001111101110000000101;
	Weight[6] = 121'b1111111100011011101111100010111100100000000000000000001111111011110001110001110011101111000011101101100000010000001011111;
	Weight[7] = 121'b1110000101011010011100010110111111000011000100001100000100011001010111001100011010111000010011100001001010001011001001111;
	Weight[8] = 121'b1010010100110100111111000011101111000110101100011100011000110101001001010001101111001110001110010110001110000000100101001;
	Weight[9] = 121'b0110000000010000000110100101101000110001001100110000110111110101100011101101000010101000100000011100000001111010001101111;
	Weight[10] = 121'b0001101001111000001100000011100010010011111110011011111111100000101111000001000110101001101010000001001011001101100011011;
	Weight[11] = 121'b0000011001010001110100100000111110000001010100000000110110101001011111101011101111001101111100000010100110100010001100101;
	Weight[12] = 121'b1101000101110111000000000101110001101110111001100000110011010011111011101111100010110011101110001000011000010110101000011;
	Weight[13] = 121'b0011110110101110011100000010011011000011000100011110000010011111001000110000000001100000000010100100000110110001010001000;
	Weight[14] = 121'b1101111000000101110011111110110000000001100011000110010001111101000010011111101010000001100000101000111010100110000000001;
	Weight[15] = 121'b0101010011110111110101110011110100110001110000000001110000001111010110000000011111111001101111110010111011101100010110101;
	Weight[16] = 121'b0100000001011101110000011101101011101011110011100111100110101101010100100000100000001101100100000000111010000110111111001;
	Weight[17] = 121'b0011011010001000010011000001000111000011111110000100001010110000000001111100010001010000111111110001000000101101000000000;
	Weight[18] = 121'b0110110111001110001101000011101000001001110101110001111011100111100111000110001110001000011101101000101100011110001010011;
	Weight[19] = 121'b0100101010101100001110100011011010001100110100011001000111110111001011101000010100010000100001100110000000110100000010000;
	Weight[20] = 121'b0010110101100000000000000111111110100111000101110000101011111010000001111000110000001101110000110111111110011111011111101;
	Weight[21] = 121'b0101011010000100100001110000111010000111111100010100001001101000010001010000010100111101000001000110000000100100011110111;
	Weight[22] = 121'b0011110110110111111010011001000011000000001010000010101000111111111111111101110110011100110000001110001010001010001000001;
	Weight[23] = 121'b0010001110001101000010010001110000000000111010001101001111010111011100001000001000100000101110000000111100000101111001001;
	Weight[24] = 121'b0000001100000010110100000000110010000111111010010001100000001100011110110001111111010011110001010111001101110100111111101;
	Weight[25] = 121'b1100000110100000000001000000000011011111111011001111111111110000110110001101100101000010100100000001011000101110111111011;
	Weight[26] = 121'b0000000000110111100001011100100001111011010011011100001011110001010101001100111100010110110110110001100000000011011111011;
	Weight[27] = 121'b1010110110100000000100011110100011111011000001111111100010000111001000001100000000101000100000000010111101010101111011100;
	Weight[28] = 121'b0100100100100110000100000100011111101111111011111001011100000000110000011001110001111010010011110111100011110111000000101;
	Weight[29] = 121'b0001110010000100001000000000100010000001110000011010011001111100001011111000100000010110000000000011001000111101010101110;
	Weight[30] = 121'b0100000000000010000100101100001101001001111101111011111011110101010000010001010001000001000110001111011011110111101000111;
	Weight[31] = 121'b1110100010011000000010000001011001000110101000000101111100101000101001011000010000100001100001100010000110000101010110110;
	Weight[32] = 121'b1000001100011101110101111011110001011100010111110100101010001100000000011000010001101100100011111110000000100110100001101;
	Weight[33] = 121'b1111010100010010010111010010011000111100000110111000100011100101110111101111101100110000110101010000101000010000110010000;
	Weight[34] = 121'b0001001010111000001111000000111000000110001110001100111010011100011001000000001010010001000110100000101111100101101011001;
	Weight[35] = 121'b0100111111111001000111100101101011101001111000101100001110011000011110001110001010001000111101001101101111011011011010100;
	Weight[36] = 121'b1101100101010111110001010100100010001010000011000000110001100000111101110011000101111111100111011001000000001100000000001;
	Weight[37] = 121'b0011000001110111100000111011000000100011000101000100001110010001010011010101100000100100010111110101111111111001011001111;
	Weight[38] = 121'b0001000001000000011000010100001100001110001111100111011000001100110000010001010011101111101110111110001000100110000000000;
	Weight[39] = 121'b1101000100000000011100110000001101111100111000011001110100011111011000010000001001110010001001110101000111111010010000001;
	Weight[40] = 121'b1010011010001000001111110110110001010011101001000010000000111111001010101010010000011000000000100011111110100111111110100;
	Weight[41] = 121'b1101001110100110011100101110101110111111000110000100001000001110001110010110101111010000111111000001010001000001111110001;
	Weight[42] = 121'b0010001110000101010010101110110010010110000110110110101000011100001100001001111100001110011111110000111010100011111001001;
	Weight[43] = 121'b1001101101100110111001010000010001111101100011100011001100011100001000110000000110011111011101010110111011101011000000011;
	Weight[44] = 121'b1110010000011001001111100000100110000101010010011011000000111110000001011000111001100001110100010110010101011101110100011;
	Weight[45] = 121'b0000110001011111101001011011100101011100100001100001001000111100010000110001111101001111100011111101100111111111111011110;
	Weight[46] = 121'b0011111110101011110010011100000001111101011111111001110101000101100011011011011000110100000010000001010111000010011101000;
	Weight[47] = 121'b0111001111101001101110011110011000100011110011011000110011100001100111000111010011111001100111110000100011001110100101000;
	Weight[48] = 121'b1111100001011001111110010101110001000000111000001100011011111001110110101100111100011011010111000001111000000001000000010;
	Weight[49] = 121'b1100011010101001111111000000100000010010100101110100000000101000001000111001000010011110010010011111100011000000100000001;
	Weight[50] = 121'b0110111011011111110011100001110011110101110001000011110100110000001011000001001100111100000111011101011010111111000100110;
	Weight[51] = 121'b0010010110001111111110110111101100111100000100000000000000000000010000010011111111111011111111011111111001011000011101010;
	Weight[52] = 121'b0100100000100100000000001011100000011111110001010011001000000101000101111000111010010101010000001110100010001001111101110;
	Weight[53] = 121'b0111101101101111111001110001101000101110000001000000010111100011100001000011010100001100101000110100100101010001101111111;
	Weight[54] = 121'b1000100010111000101000011110111110111000101100110000000111110001001001011100000001001110000000011100010011010101000110000;
	Weight[55] = 121'b1111111111110111110010011110001110011101000001111000110001010011100011100011100011100100110011101010001000101100011001010;
	Weight[56] = 121'b0110100000110101110111100000001110001110111100111000000110010001001000100111100100011100010111110111101111110101011000111;
	Weight[57] = 121'b1111111011110100111001010001001000110011000000001011000011111011111011101101100101101100110110000011000000000011000110100;
	Weight[58] = 121'b0001101001110111000011111111111111000011101010000001011110100010000000000111011000000011110111100101111111101100011111101;
	Weight[59] = 121'b1101110110011110011100001101011001001101110001100011101100000100011100110101011001100011111111010011010100010011011111010;
		
	
	
	//Loading weight [10,64] : [output,input]
	Weight_out[0] = 60'b011001010011110001000001010001000011100010000101101001011110;
	Weight_out[1] = 60'b011000010001011010101100101000111010111000111000010001000101;
	Weight_out[2] = 60'b011000100001101100000010111111000110111000010100111110001111;
	Weight_out[3] = 60'b000110010000001110001001101001000001010111110101111011010111;
	Weight_out[4] = 60'b100010011100011001110011001001110100100110111001001000100100;
	Weight_out[5] = 60'b000100011010000001001111110011110011000011100100100101111010;
	Weight_out[6] = 60'b000100111000010001000011100010001111100010001111110001010100;
	Weight_out[7] = 60'b011010010010011010000111011110111100000011010011001011000011;
	Weight_out[8] = 60'b110101001110111010001000100010011011000101010100110000010000;
	Weight_out[9] = 60'b101000000100110110111101110101010010000010101101100011010000;
 
	
	
	/*	//****** Prueba con red del paper ******
	//Loading weight [60,121] : [output,input] without BatchNormalization Accuracy of 84.4% / implementation Accuracy of 82%
	Weight[0] = 121'b1111111100110011111100000011111101111111111011100111111011001011110001110011101111111111111111111110111111001011111111111;
	Weight[1] = 121'b1101100001100010000010000000001110000000000100000000000011111000001011000010001111001000000000011010000000111011000001100;
	Weight[2] = 121'b0010011010010000001111000000001110000000000110110000000011000000011000111000000001010000000000000000000000110000000011100;
	Weight[3] = 121'b1110111111011010110001100001000000000010000000010100000000101111010000110000010111110000000001100000000000000100000000111;
	Weight[4] = 121'b1011110111011111100000101100000000000000000000000010000000001100001000110001100001000011000000001111110000010111100000101;
	Weight[5] = 121'b1000000000100000000001100000000000000000000000000000000100000000001000000000010000000000100000000001100000000011000000011;
	Weight[6] = 121'b0000000000010000000000100000000000000000000000000000000000000000001000000000000000000000100000000001100000000011000000000;
	Weight[7] = 121'b0111111111111111111010100111110000011111111000111111000001111111100111111111010011111101110111110111001011100100001100011;
	Weight[8] = 121'b1011011000000000000000100000000000000000000000000000000100000000000000010000000000000001000000000010000000001111000011011;
	Weight[9] = 121'b0011100011010000000011110000111101101100111011111001110111100001110011000011000110000000001100100000001010001111110010010;
	Weight[10] = 121'b0000000000110000000000000000000011000000000011100000000110000000000000000000000000000000100000000001000000100010000011101;
	Weight[11] = 121'b1101101110111111100001111100000001100000000000000010000000000000001000000000100000000110011000001101111100000001111100000;
	Weight[12] = 121'b0010100110010000000001100000000000000000000000000000011000000000110000000000110000000000100000000010000000000110000000001;
	Weight[13] = 121'b0010001111000101011110011100000010110000000100000000000000000011001000000010010011100100110111001101111100010011111000000;
	Weight[14] = 121'b1000011000110000010000100000001001111110001011111000100111000000110000011000000110110000000001100000000001000000001110100;
	Weight[15] = 121'b1011110000100001100001000110000000010000000000010000000000100000000001000110000000010000000010010000000100000010010000010;
	Weight[16] = 121'b1100000010000000000100000001100010000000000100000100111000111000000011100010101111001000110110010000000000100000000000110;
	Weight[17] = 121'b0110000000100100000011101110011110000000001100000000001000011000001000100000010000000000111100011101111000111111100001111;
	Weight[18] = 121'b0001111110001111100000010001000101101100010010111001110111100011111011001110010010011100110001110001000000010011001011000;
	Weight[19] = 121'b0000000000110000000001000000000000000000000000000000000100000000001000000000000000000000000000000011000000000010000000001;
	Weight[20] = 121'b0001001111001000010001110000000101100001000000001110000000010000001000000010011000000000011011000100110000001000000000011;
	Weight[21] = 121'b1100000000110000000001100000001110001000000100100000100010000000001000000000100000000000000000000000000000111010000011110;
	Weight[22] = 121'b0100100100010000000001100000000000000000000000000000001000000000010000000000100000000000000000000000000000000000000000000;
	Weight[23] = 121'b0100011001001001000011110000000010000010000010000000001100000000101100000001001100000010000100000011010100000011101000000;
	Weight[24] = 121'b1000000000110000000001000000000001110110011011100000110110000000000000000000010000000000000000000011000011001110011111011;
	Weight[25] = 121'b0000000001100100000001100000000110000000011100000000111000000000001000000000001000000000110000001110000000011011000000000;
	Weight[26] = 121'b1011111111001111010011111110111011111110110100111111001110111111111011111111110111111111101111111011001101111111111111111;
	Weight[27] = 121'b1000100001000111100000011100000100000000000010000000000000000000011100000011010000000110101110001110111110001110011100000;
	Weight[28] = 121'b1100000000010000000000100000000010000000001100100000011110000000110110000000010000000000000000000001000000000100000001101;
	Weight[29] = 121'b1001000001000111000000101110010000010001100000000110001000000000001100000110001000000110011110011000011110000001111100000;
	Weight[30] = 121'b0000000000010010110000011111110001101111110001110111110001111111110011111111101011110011001011111010001101100011111110000;
	Weight[31] = 121'b1101100111010000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
	Weight[32] = 121'b0100000000010000000001000000000000000000000000000000000100000000001000000000000000000000000000000000100000000000111000000;
	Weight[33] = 121'b0110100000100000100000000000100000000011000000000110000000011000000000010000000001100000000011000000000101000010000000000;
	Weight[34] = 121'b0100000001001001010011000101011110101101011100111011110011110111001001101000000000000100010101000000010111111000000000100;
	Weight[35] = 121'b1010000001010000000001100000000011000000000100000000000100000000000000000000010000000000100000000011100000000101000000001;
	Weight[36] = 121'b1000000000000000000001010000000000000000000000000000000000000000000000000000001000000000011000000010111100000110111100011;
	Weight[37] = 121'b0000000011100000000000000001100000000001001000100110011000001000000010011000000001110000000011000000000000000001001100000;
	Weight[38] = 121'b0010111110010011110000000000000000000000000100000000000000000000011000000000110000000000100000000010000000000010000000000;
	Weight[39] = 121'b1011000111010000101111001001011110111010010110111010011100011110100011111010000101001000000011101000000100100011000101011;
	Weight[40] = 121'b1010000000101100000000011110000100111111111110010111011111000000011100011100010110100000000100000000000111000000101110011;
	Weight[41] = 121'b0010011000000000101001001110111110001101011100111101011011101000000010110000000110000110001111110100000101111010000000010;
	Weight[42] = 121'b0110111111000111111100001010000010000000000100000000111010000001110011000011101110001110001100011100110000010010000000000;
	Weight[43] = 121'b1011111111011101011100111001111111111101101010101111100101101010111001111010010001011010000001010000000011000001100001100;
	Weight[44] = 121'b1100010000011101110000101111110101100011110100100110110000011111011110010110111010001110101110110001001011010100000000001;
	Weight[45] = 121'b1111101111010101010111000110100010000100001100111000110001110011100001101011010111101110000111100101101011100010000000010;
	Weight[46] = 121'b1100101000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000100000000000000000000;
	Weight[47] = 121'b0000000111100010011111001000110111000011001000001110000100010000100100000010000000000110010111000000001100000000101000100;
	Weight[48] = 121'b1001000011101000000111001110011000001001110010000011100101000111001001001011000001000000001110000000011100000111001000000;
	Weight[49] = 121'b1011011011011011000000000000000010000000000100000000001000000000111000000001101100000011011000001111000000010010000000111;
	Weight[50] = 121'b0100000001000000000000100001100001000011000000000110001110000000001100010000011000000001100010000010000011001100000000011;
	Weight[51] = 121'b1111101110101111110110111110111111100101000000110001110101110010111101100110100111100111001111111011101010000100000000001;
	Weight[52] = 121'b1111110001010000000001000101010000011111000000111000000000100110000000100100000000011001000001010010000111110100001111111;
	Weight[53] = 121'b1100000100111001100001111111111100110111111110111111101101110011001111000111010100011100111011010101111111000011110111111;
	Weight[54] = 121'b1000000000000010000000101110001111011001110100000111000000000010000100000100000000000000000010011001011100100010100000111;
	Weight[55] = 121'b1011000111100000000011000001111000000111101000111100100000101010110111000100000011001000001011000000000111010000000011110;
	Weight[56] = 121'b1010000001101110000001000000000000000000000010000000000110000000011000000000000000000001100000000101000000001111000000111;
	Weight[57] = 121'b0100000010000000001011000001101010011111000011110000010111110001100000000011000100100010000101000000001011100110001011001;
	Weight[58] = 121'b1011111100100110110011110000000000100000000000000000000110000000001100000011111011000111100000000110000000000101000000011;
	Weight[59] = 121'b1110000010100000000011000000000000000000000000000000000100000000001000000000000000000000000000000001100000000011100000000;
	

	Weight_out[0] = 60'b111111111111111111011111100010111100111100100111011111110111;
	Weight_out[1] = 60'b110101110001111111100110111111011101110011111011111010111111;
	Weight_out[2] = 60'b100000010000000100000000001100100100010000000000000110000000;
	Weight_out[3] = 60'b100000010100001000010000001011000100010000011000000011001000;
	Weight_out[4] = 60'b011011111111111001111111111111111011101100110011011100000111;
	Weight_out[5] = 60'b111101111011111111010111111111010101111111100111010011111111;
	Weight_out[6] = 60'b111111111011111111111111111111011101111110110111011110111111;
	Weight_out[7] = 60'b111011101111111111110111111111111101111110110011111011110111;
	Weight_out[8] = 60'b100100000000000100000000001000100110100101011100000010010100;
	Weight_out[9] = 60'b111001111011111101110111111111111111111000100011011010111011;   */

	/*	//****** Prueba con red del paper ******
	//Loading weight [48,121] : [output,input] with BatchNormalization Accuracy of 94.3% / implementation Accuracy of %
	Weight[0] = 121'b0011011110010111111111000111110100110100000000000000010001110001111010100101010011111111010111111110010000010011001000011;
	Weight[1] = 121'b0111111001100111111011100010010000001010111111000110111000000000011000010011111111110001111111111010100000110100000001001;
	Weight[2] = 121'b0111101000110110101101011000111011001011101110001110001100111100000100001000101100110001011110000010111000001111110001110;
	Weight[3] = 121'b1010110101000011000000101111000011111111000011110001001010000110010000011000100001111010100111001010010001011110011111101;
	Weight[4] = 121'b1111011101001001111111100000011010100000010110010110110100001100100001010000000001111110100111111000100011100010000000011;
	Weight[5] = 121'b0110000111001000010111000000001111000010011101001100100010011000001000110000000110110000100011100011000100100000001000100;
	Weight[6] = 121'b0010110010111101100010100010000100111000010001111001110011101111101100111000000000111001011000010011111100110000111010101;
	Weight[7] = 121'b1000000101011001110001111100010010101001100010101111000110000000001100001110110000011000010011110000011111011101111111100;
	Weight[8] = 121'b1100010100011111010010010001110001000101111000101101110110101011101111100010110110000011011111000010001100100010101010000;
	Weight[9] = 121'b1110001001101001000000000001110010000101111110001000000100111100010100101100011000011011111001100010101110000011011111111;
	Weight[10] = 121'b0100000000100000001100011010010110111110010111011010000100110111000111001110011000100100110001000010100110111011110000000;
	Weight[11] = 121'b0111100000111110100011100111100100000111111101000000011100000001111001100010100111100011011101111100111111111010001000011;
	Weight[12] = 121'b0101010010000101111101100010100000100010010000001100110001010000101011000111001111110111101101111101000111010100100100100;
	Weight[13] = 121'b1001010000001111110010110111111001110010000111001001011100111101011000000010100000011111110111010101111111101100111111011;
	Weight[14] = 121'b0111010110001000101100001001111010000110000000101101000000111111001000111000010011000000100011000100000100000111000111100;
	Weight[15] = 121'b0110000110010100000000101011100010000010100101011110000110011101100000011000110010100001111000110010001010100010100001100;
	Weight[16] = 121'b0100100100001000001000111100111000101001000000111011100011110111010011101100110000010001000000100011010001010001110111101;
	Weight[17] = 121'b1001010000001111100000010011100101001011001111100101100000001100000100110000010011001100010010111110100111110110010100000;
	Weight[18] = 121'b0110010110111110001011011001011110100010101100011100001011110001100101000111011000001111010111010100000111111001011011110;
	Weight[19] = 121'b0001000011111111110000001000001000100001000110001000100101110001111111101111101111111000111111001110000001001010000000010;
	Weight[20] = 121'b1011101000111010110011000111101000011011100101110010111110111111111100000111010110001110001101111101001010111011111100111;
	Weight[21] = 121'b0000000010101000001101001100000110011100101100011000100111010010010101011110111100011001101011111100111111011111010000001;
	Weight[22] = 121'b1111111010011000011010011001111001011101110100000011000000001101001000110001111011101001111111011110010000001001111010101;
	Weight[23] = 121'b1101111011010110000011110000011001000110000010011001000001111110010111111000001011000010100000111100010000111001111110110;
	Weight[24] = 121'b1001100011000101010110110111100110101000011110110001110100111100110001100001000001010110100010100001100011111111101101100;
	Weight[25] = 121'b1110000011000111101110000010101000100110001011101110000010001011011100010001111011111110111111111110110100001011000001010;
	Weight[26] = 121'b1011111111000011111100011000110001001110000100000000000010011101110111111111100011100110011101010001100001010010110010000;
	Weight[27] = 121'b0000001111100001101011110000110110000100000010010001011010110111110011111010111100111111010100011110000000111101111100000;
	Weight[28] = 121'b1011101100101000000000100000100011000111111110101000111011110000000010000100010011100001000000010100110100001011111111111;
	Weight[29] = 121'b0100010000001111101011010111110010101011010000010001100100000000000110000100111101110010111101111111101100111011011111110;
	Weight[30] = 121'b1000000110111000111111000000011111011100111110011000001111111101000100011001010001000011000000111001000011010111000000011;
	Weight[31] = 121'b0001010100110010111110110011101010100000111100001100011110011000011111001100111110011000110111001101100100000011100001110;
	Weight[32] = 121'b0110111000001000111110000111101110001110000110110100001011000010001100000000011100011011011001111111101101111001011001110;
	Weight[33] = 121'b1110111110110110001110001100000010111100000001011000010001010011100000110000010011110001100111111101000111010011100010010;
	Weight[34] = 121'b1110110011111000000000000000111011001011001101011000111001111001110010101001101111010111111100000001001110010000101111111;
	Weight[35] = 121'b1100111110010001001110000000111110000110001100001111010101010001101011000011001110010000001111010001001010000010100000001;
	Weight[36] = 121'b1111110010001101111100000101110001000100111001000001100000011000010110110000111110011000101011100011011111101111011011101;
	Weight[37] = 121'b0100111111001111000010101100000011110110001001000100000000011010001010110111011000011110111100110011111111100000111110101;
	Weight[38] = 121'b1011110001000011010010000011001010110000101010001010000011110111111011011111010001011111001100000000001100001110110100011;
	Weight[39] = 121'b1100000100011100100000100011111011000111111010010011110010101110001100011000001001010000011000000000010010000111111111111;
	Weight[40] = 121'b1001010101100001111001100000011101110111111001101001111000100010100001000000100011000011011010010000010110100010000110011;
	Weight[41] = 121'b1101000010110111110010101111110101011000001101111101000001011010010000111101011010001101100100011101101110111011011011011;
	Weight[42] = 121'b0101011110100000111111000011110011101110000000011000000011110111001001100100010011001000011001100000100011111110001111110;
	Weight[43] = 121'b0011000001110000100010110110010111000110111100001100011000101100010100011000000111111001100110000110001111000101001010000;
	Weight[44] = 121'b1001000000010011111000011010110000100001100000000010000011111010011111101000110110011101101100010101101001101100010000001;
	Weight[45] = 121'b0001101010000111100001010100011100101001100000010011111111100101101110000011100010011100101110100010111001100110011101110;
	Weight[46] = 121'b0101100111111001000000110011010000001011100100110001100011010011100111101101100011011000110101001110100101011011101001110;
	Weight[47] = 121'b0110100100010000000101011111000011110111000011000111000110101001111100010101010100000111100000000111000100000101111111101;




	Weight_out[0] = 48'b101000001101101001110000100000011010100010100110;
	Weight_out[1] = 48'b011011000000110101000111010000001010000010001101;
	Weight_out[2] = 48'b110100000001010001010111111101110010101010001001;
	Weight_out[3] = 48'b011000110100110001111011110001010000110100001001;
	Weight_out[4] = 48'b101001100011101110010101100101100001001000011000;
	Weight_out[5] = 48'b111001000101010010100100110110111011000001110000;
	Weight_out[6] = 48'b101011100000101001110001101100010101001000100100;
	Weight_out[7] = 48'b000100110010100111100010001011000000001110110101;
	Weight_out[8] = 48'b000010111001001101001000110100110111100111111000;
	Weight_out[9] = 48'b001000101100011110001001100110001001000100110011;


    
	scaling[0] = 4'd2;
	scaling[1] = 4'd2;
	scaling[2] = 4'd2;
	scaling[3] = 4'd2;
	scaling[4] = 4'd2;
	scaling[5] = 4'd1;
	scaling[6] = 4'd2;
	scaling[7] = 4'd2;
	scaling[8] = 4'd2;
	scaling[9] = 4'd2;
	scaling[10] = 4'd2;
	scaling[11] = 4'd2;
	scaling[12] = 4'd2;
	scaling[13] = 4'd2;
	scaling[14] = 4'd2;
	scaling[15] = 4'd2;
	scaling[16] = 4'd2;
	scaling[17] = 4'd2;
	scaling[18] = 4'd2;
	scaling[19] = 4'd2;
	scaling[20] = 4'd2;
	scaling[21] = 4'd2;
	scaling[22] = 4'd2;
	scaling[23] = 4'd2;
	scaling[24] = 4'd2;
	scaling[25] = 4'd2;
	scaling[26] = 4'd2;
	scaling[27] = 4'd2;
	scaling[28] = 4'd2;
	scaling[29] = 4'd2;
	scaling[30] = 4'd2;
	scaling[31] = 4'd2;
	scaling[32] = 4'd2;
	scaling[33] = 4'd3;
	scaling[34] = 4'd2;
	scaling[35] = 4'd2;
	scaling[36] = 4'd2;
	scaling[37] = 4'd2;
	scaling[38] = 4'd3;
	scaling[39] = 4'd2;
	scaling[40] = 4'd2;
	scaling[41] = 4'd2;
	scaling[42] = 4'd2;
	scaling[43] = 4'd2;
	scaling[44] = 4'd2;
	scaling[45] = 4'd2;
	scaling[46] = 4'd2;
	scaling[47] = 4'd2;



	offset[0] = 4'b0;
	offset[1] = 4'b10;
	offset[2] = 4'b10;
	offset[3] = 4'b10;
	offset[4] = 4'b10;
	offset[5] = 4'b110;
	offset[6] = 4'b10;
	offset[7] = 4'b10;
	offset[8] = 4'b1110;
	offset[9] = 4'b1110;
	offset[10] = 4'b0;
	offset[11] = 4'b0;
	offset[12] = 4'b0;
	offset[13] = 4'b0;
	offset[14] = 4'b0;
	offset[15] = 4'b10;
	offset[16] = 4'b10;
	offset[17] = 4'b0;
	offset[18] = 4'b10;
	offset[19] = 4'b100;
	offset[20] = 4'b1011;
	offset[21] = 4'b0;
	offset[22] = 4'b1110;
	offset[23] = 4'b10;
	offset[24] = 4'b10;
	offset[25] = 4'b1110;
	offset[26] = 4'b0;
	offset[27] = 4'b10;
	offset[28] = 4'b1010;
	offset[29] = 4'b10;
	offset[30] = 4'b101;
	offset[31] = 4'b10;
	offset[32] = 4'b110;
	offset[33] = 4'b11;
	offset[34] = 4'b10;
	offset[35] = 4'b100;
	offset[36] = 4'b0;
	offset[37] = 4'b101;
	offset[38] = 4'b0;
	offset[39] = 4'b1110;
	offset[40] = 4'b1000;
	offset[41] = 4'b1110;
	offset[42] = 4'b1110;
	offset[43] = 4'b1110;
	offset[44] = 4'b10;
	offset[45] = 4'b101;
	offset[46] = 4'b1110;
	offset[47] = 4'b1000;   */
	
    
	   
  end
  
  
  //********** Using Generate **********
  
  localparam size_weight = 1;
  
  genvar i;
  generate
  
   // First Hidden Layer 128 neuron
  for(i=0;i<number_output1;i=i+1)begin
    neuron#(size_word,number_image,size_weight) h1(
        .Image(Image),
        .Weight(Weight[i]),
        .out(out_aux[(2*size_word)*(i+1)-1:2*size_word*i])
    );
  end 
  
 
  
   // Ouput Layer 10
  for(i=0;i<number_out;i=i+1)begin
    neuron_out#(2*size_word,number_output1,size_weight) out(
        .Image(out_aux),
        .Weight(Weight_out[i]),
        .out(out_aux_out[(4*size_word)*(i+1)-1:4*size_word*i])
    );
  end 

  
  
  wire signed [31:0] out_test [9:0];
   
  for(i=0; i<10; i=i+1)begin
        assign out_test[i] = out_aux_out[32*(i+1)-1:32*i];
  end 
  


 endgenerate 
 //*****************************************************
    
  //*********** Prediction Function **********
  
  reg signed [31:0] maximux;
  reg [3:0] prediction;
  integer j;
  always@(*)begin
    maximux = out_test[0];
    prediction = 0;
    for(j=1;j<10;j=j+1)begin
        if(out_test[j] > maximux) begin
            maximux = out_test[j];
            prediction = j;
        end
    end
  
  end
 
  assign regr_0 = prediction;
  //*******************************************************************************

endmodule